** sch_path: /home/herman/github/KrzysztofHerman/IHP-Open-DesignLib/ts_pr_May2024/design_data/xschem/transmission_gate_v1.sch
.subckt ESD-2kv vdd inout_1 inout_2 vss en
*.PININFO inout_1:B inout_2:B en:I vdd:B vss:B
M1 inout_2 net1 inout_1 sub sg13_lv_nmos L=0.130u W=5.0u ng=5 m=1
M2 inout_1 en inout_2 nwell sg13_lv_pmos L=0.130u W=5.0u ng=5 m=1
R1 vss sub ptap1 l=780n w=780n
R2 vdd nwell ntap1 l=780n w=780n
M3 net1 en vss sub sg13_lv_nmos L=0.130u W=0.740u ng=1 m=1
M4 net1 en vdd nwell sg13_lv_pmos L=0.130u W=1.120u ng=1 m=1
D1 sub en dantenna l=780n w=780n
D2 en nwell dpantenna l=780n w=780n
.ends
.end
