** sch_path: /home/herman/github/KrzysztofHerman/IHP-Open-DesignLib/ts_pr_May2024/design_data/xschem/resistors_tb.sch
**.subckt resistors_tb
Vres Vcc GND 1.5
Vsil Vcc net2 0
.save i(vsil)
Vppd net4 GND 0
.save i(vppd)
Vrh Vcc net3 0
.save i(vrh)
Vptap net5 GND 0
.save i(vptap)
Vntap Vcc net1 0
.save i(vntap)
x1 Vcc net1 net3 Vcc net2 net5 GND net4 GND GND resistors
**** begin user architecture code

.lib /home/herman/github/KrzysztofHerman/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ



.param temp=27
.control
save all
op
echo Silicide resisotr value:
print Vcc/I(Vsil)
echo Unsilicide poly resisotr value:
print Vcc/I(Vppd)
echo High poly resisotr value:
print Vcc/I(Vrh)
reset
dc temp -40 125 1
write dc_res_temp.raw
wrdata dc_res_temp.csv I(Vsil) I(Vppd) I(Vrh)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  resistors.sym # of pins=10
** sym_path: /home/herman/github/KrzysztofHerman/IHP-Open-DesignLib/ts_pr_May2024/design_data/xschem/resistors.sym
** sch_path: /home/herman/github/KrzysztofHerman/IHP-Open-DesignLib/ts_pr_May2024/design_data/xschem/resistors.sch
.subckt resistors rppd_p ntap1_p rhigh_p ptap1_p rsil_p ptap1_n rhigh_n rppd_n rsil_n ntap1_n
*.iopin ntap1_p
*.iopin ptap1_p
*.iopin rsil_p
*.iopin rppd_p
*.iopin rhigh_p
*.iopin ntap1_n
*.iopin ptap1_n
*.iopin rsil_n
*.iopin rppd_n
*.iopin rhigh_n
XR2 rppd_n rppd_p rppd w=0.5e-6 l=2.5e-6 m=1 b=0
XR3 rhigh_n rhigh_p rhigh w=0.5e-6 l=2.0e-6 m=1 b=0
XR1 rsil_n rsil_p rsil w=0.5e-5 l=0.5e-5 m=1 b=0
XR4 ptap1_n ptap1_p ptap1
XR5 ntap1_n ntap1_p ntap1
.ends

.GLOBAL GND
.end
