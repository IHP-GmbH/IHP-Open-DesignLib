// Licensed to the Apache Software Foundation (ASF) under one
// or more contributor license agreements.  See the NOTICE file
// distributed with this work for additional information
// regarding copyright ownership.  The ASF licenses this file
// to you under the Apache License, Version 2.0 (the
// "License"); you may not use this file except in compliance
// with the License.  You may obtain a copy of the License at

//   http://www.apache.org/licenses/LICENSE-2.0

// Unless required by applicable law or agreed to in writing,
// software distributed under the License is distributed on an
// "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY
// KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations
// under the License.    

`define SIZE 1600

module shreg(
    clk,
    rst,
    shreg_enable,
    shreg_in,
    shreg_out
);

input wire clk;
input wire rst;
input wire shreg_enable;
input wire shreg_in;
output wire shreg_out;

reg [`SIZE-1:0] storage; 

always @(posedge clk) begin
    if(rst == 1'b0) 
        storage <= {`SIZE{1'b0}};
    else if (shreg_enable == 1'b1)
        storage <= {storage[`SIZE-2:0], shreg_in};
    else
        storage <= storage;
end

assign shreg_out = storage[`SIZE-1];

endmodule
