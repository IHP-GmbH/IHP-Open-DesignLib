** sch_path: /home/herman/github/KrzysztofHerman/IHP-Open-DesignLib/ts_pr_May2024/design_data/xschem/transmission_gate_tb.sch
**.subckt transmission_gate_tb
Vpow net1 GND 1.2
Vp net1 net2 0
.save i(vp)
x1 net2 V_in V_out GND en_in transmission_gate_v1
Vin V_in GND dc=0 ac=1 sin(0, 200m, 20meg, 0, 0)
Ven en_in GND pulse(0 1.2 0 1p 1p 50n 100n)
C1 V_out GND 10p m=1
**** begin user architecture code

.lib /home/herman/github/KrzysztofHerman/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.include /home/herman/github/KrzysztofHerman/IHP-Open-PDK/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27
.control
pre_osdi ./psp103_nqs.osdi
save all
tran 1p 120n
write tran_res_temp.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  transmission_gate_v1.sym # of pins=5
** sym_path: /home/herman/github/KrzysztofHerman/IHP-Open-DesignLib/ts_pr_May2024/design_data/xschem/transmission_gate_v1.sym
** sch_path: /home/herman/github/KrzysztofHerman/IHP-Open-DesignLib/ts_pr_May2024/design_data/xschem/transmission_gate_v1.sch
.subckt transmission_gate_v1 vdd inout_1 inout_2 vss en
*.iopin inout_1
*.iopin inout_2
*.ipin en
*.iopin vdd
*.iopin vss
x1 en VDD VSS net1 sg13g2_inv_1
XM1 inout_2 net1 inout_1 vss sg13_lv_nmos W=5.0u L=0.130u ng=1 m=1
XM2 inout_1 en inout_2 vdd sg13_lv_pmos W=5.0u L=0.130u ng=1 m=1
.ends

.GLOBAL GND
.end
