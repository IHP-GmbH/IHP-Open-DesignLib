* Extracted by KLayout with SG13G2 LVS runset on : 25/04/2024 17:23

* cell TOP
.SUBCKT TOP
.ENDS TOP
