module riscv (clk,
    memread,
    memwrite,
    reset,
    suspend,
    aluout,
    instr,
    pc,
    readdata,
    writedata);
 input clk;
 output memread;
 output memwrite;
 input reset;
 output suspend;
 output [31:0] aluout;
 input [31:0] instr;
 output [31:0] pc;
 input [31:0] readdata;
 output [31:0] writedata;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire net170;
 wire net169;
 wire net168;
 wire net167;
 wire net166;
 wire net165;
 wire net164;
 wire net163;
 wire net162;
 wire net161;
 wire net160;
 wire net159;
 wire net158;
 wire net157;
 wire net156;
 wire net155;
 wire net154;
 wire net153;
 wire net152;
 wire net151;
 wire net150;
 wire net149;
 wire net148;
 wire net147;
 wire net146;
 wire net145;
 wire net144;
 wire net143;
 wire net142;
 wire net141;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire net104;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire net103;
 wire _02089_;
 wire net102;
 wire _02091_;
 wire _02092_;
 wire net101;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire net100;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire net99;
 wire net98;
 wire net97;
 wire _02115_;
 wire net96;
 wire _02117_;
 wire net95;
 wire _02119_;
 wire net94;
 wire _02121_;
 wire _02122_;
 wire net93;
 wire net92;
 wire net91;
 wire _02126_;
 wire net90;
 wire _02128_;
 wire net89;
 wire _02130_;
 wire net88;
 wire _02132_;
 wire net87;
 wire _02134_;
 wire net86;
 wire _02136_;
 wire net85;
 wire net84;
 wire _02139_;
 wire net83;
 wire _02141_;
 wire _02142_;
 wire net82;
 wire _02144_;
 wire net81;
 wire net80;
 wire _02147_;
 wire _02148_;
 wire net79;
 wire _02150_;
 wire net78;
 wire _02152_;
 wire _02153_;
 wire net77;
 wire _02155_;
 wire _02156_;
 wire net76;
 wire _02158_;
 wire net75;
 wire _02160_;
 wire net74;
 wire _02162_;
 wire net73;
 wire _02164_;
 wire net72;
 wire _02166_;
 wire net71;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire net70;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire net69;
 wire net68;
 wire net67;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire net66;
 wire _02187_;
 wire _02188_;
 wire net65;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire net64;
 wire _02199_;
 wire _02200_;
 wire net63;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire net62;
 wire net61;
 wire net60;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire net59;
 wire _02225_;
 wire _02226_;
 wire net58;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire net57;
 wire _02237_;
 wire _02238_;
 wire net56;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire _02255_;
 wire _02256_;
 wire net51;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire net50;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire net49;
 wire _02269_;
 wire _02270_;
 wire net48;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire net47;
 wire net46;
 wire _02293_;
 wire _02294_;
 wire net45;
 wire net44;
 wire net43;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire net42;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire net41;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire net40;
 wire net39;
 wire net38;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire net37;
 wire _02342_;
 wire _02343_;
 wire net36;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire net35;
 wire _02354_;
 wire _02355_;
 wire net34;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire net33;
 wire net32;
 wire net31;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire net30;
 wire _02380_;
 wire _02381_;
 wire net29;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire net28;
 wire _02392_;
 wire _02393_;
 wire net27;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire net26;
 wire _02407_;
 wire _02408_;
 wire net25;
 wire net24;
 wire net23;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire net22;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire net21;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire net20;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire net19;
 wire net18;
 wire net17;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire net16;
 wire _02457_;
 wire _02458_;
 wire net15;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire net14;
 wire _02469_;
 wire _02470_;
 wire net13;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire net12;
 wire net11;
 wire net10;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire net9;
 wire _02495_;
 wire _02496_;
 wire net8;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire net7;
 wire _02507_;
 wire _02508_;
 wire net6;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire net5;
 wire net4;
 wire net3;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire net2;
 wire _02533_;
 wire _02534_;
 wire net1;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02545_;
 wire _02546_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire net1161;
 wire _02559_;
 wire net1160;
 wire _02561_;
 wire net1159;
 wire net1158;
 wire net1157;
 wire _02565_;
 wire net1156;
 wire net1155;
 wire net1154;
 wire net1153;
 wire _02570_;
 wire net1152;
 wire _02572_;
 wire net1151;
 wire net1150;
 wire net1149;
 wire _02576_;
 wire net1148;
 wire _02578_;
 wire net1147;
 wire net1146;
 wire net1145;
 wire net1144;
 wire _02583_;
 wire net1143;
 wire net1142;
 wire net1141;
 wire net1140;
 wire net1139;
 wire net1138;
 wire net1137;
 wire net1136;
 wire _02592_;
 wire _02593_;
 wire net1135;
 wire net1134;
 wire net1133;
 wire _02597_;
 wire _02598_;
 wire net1132;
 wire net1131;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire net1130;
 wire _02605_;
 wire net1129;
 wire net1128;
 wire net1127;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire net1126;
 wire net1125;
 wire net1124;
 wire _02615_;
 wire _02616_;
 wire net1123;
 wire net1122;
 wire net1121;
 wire _02620_;
 wire net1120;
 wire net1119;
 wire net1118;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire net1117;
 wire net1116;
 wire net1115;
 wire _02630_;
 wire _02631_;
 wire net1114;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire net1113;
 wire _02637_;
 wire net1112;
 wire net1111;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire net1110;
 wire net1109;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire net1108;
 wire _02649_;
 wire net1107;
 wire net1106;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire net1105;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire net1104;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire net1103;
 wire net1102;
 wire _02673_;
 wire _02674_;
 wire net1101;
 wire net1100;
 wire _02677_;
 wire net1099;
 wire net1098;
 wire net1097;
 wire net1096;
 wire net1095;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire net1094;
 wire net1093;
 wire net1092;
 wire net1091;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire net1090;
 wire _02695_;
 wire _02696_;
 wire net1089;
 wire net1088;
 wire _02699_;
 wire net1087;
 wire _02701_;
 wire _02702_;
 wire net1086;
 wire net1085;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire net1084;
 wire net1083;
 wire _02711_;
 wire _02712_;
 wire net1082;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire net1081;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire net1080;
 wire net1079;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire net1078;
 wire net1077;
 wire net1076;
 wire _02735_;
 wire net1075;
 wire _02737_;
 wire _02738_;
 wire net1074;
 wire net1073;
 wire _02741_;
 wire _02742_;
 wire net1072;
 wire net1071;
 wire _02745_;
 wire _02746_;
 wire net1070;
 wire _02748_;
 wire net1069;
 wire net1068;
 wire net1067;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire net1066;
 wire net1065;
 wire net1064;
 wire _02758_;
 wire _02759_;
 wire net1063;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire net1062;
 wire _02770_;
 wire net1061;
 wire net1060;
 wire net1059;
 wire _02774_;
 wire net1058;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire net1057;
 wire net1056;
 wire net1055;
 wire _02785_;
 wire _02786_;
 wire net1054;
 wire _02788_;
 wire _02789_;
 wire net1053;
 wire net1052;
 wire _02792_;
 wire _02793_;
 wire net1051;
 wire _02795_;
 wire net1050;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire net1049;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire net1048;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire net1047;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire net1046;
 wire _02822_;
 wire net1045;
 wire net1044;
 wire net1043;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire net1042;
 wire net1041;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire net1040;
 wire _02850_;
 wire net1039;
 wire _02852_;
 wire _02853_;
 wire net1038;
 wire _02855_;
 wire _02856_;
 wire net1037;
 wire _02858_;
 wire _02859_;
 wire net1036;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire net1035;
 wire _02867_;
 wire _02868_;
 wire net1034;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire net1033;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire net1032;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire net1031;
 wire _02900_;
 wire net1030;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire net1029;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire net1028;
 wire net1027;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire net1026;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire net1025;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire net1024;
 wire _02976_;
 wire net1023;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire net1022;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire net1021;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire net1020;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire net1019;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire net1018;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire net1017;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire net1016;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire net1015;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire net1014;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire net1013;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire net1012;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire net1011;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire net1010;
 wire net1009;
 wire net1008;
 wire _03133_;
 wire _03134_;
 wire net1007;
 wire _03136_;
 wire _03137_;
 wire net1006;
 wire _03139_;
 wire _03140_;
 wire net1005;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire net1004;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire net1003;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire net1002;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire net1001;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire net1000;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire net999;
 wire net998;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire net997;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire net996;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire net995;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire net994;
 wire _03303_;
 wire _03304_;
 wire net993;
 wire net992;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire net991;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire net990;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire net989;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire net988;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire net987;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire net986;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire net985;
 wire net984;
 wire net983;
 wire _03654_;
 wire net982;
 wire net981;
 wire net980;
 wire net979;
 wire net978;
 wire net977;
 wire net976;
 wire _03662_;
 wire net975;
 wire net974;
 wire net973;
 wire _03666_;
 wire net972;
 wire net971;
 wire net970;
 wire net969;
 wire net968;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire net967;
 wire _03676_;
 wire net966;
 wire net965;
 wire net964;
 wire _03680_;
 wire _03681_;
 wire net963;
 wire _03683_;
 wire net962;
 wire _03685_;
 wire _03686_;
 wire net961;
 wire net960;
 wire _03689_;
 wire net959;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire net958;
 wire net957;
 wire net956;
 wire _03697_;
 wire _03698_;
 wire net955;
 wire net954;
 wire _03701_;
 wire _03702_;
 wire net953;
 wire net952;
 wire _03705_;
 wire net951;
 wire _03707_;
 wire net950;
 wire net949;
 wire net948;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire net947;
 wire _03719_;
 wire net946;
 wire _03721_;
 wire net945;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire net944;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire net943;
 wire net942;
 wire net941;
 wire _03734_;
 wire _03735_;
 wire net940;
 wire _03737_;
 wire net939;
 wire net938;
 wire net937;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire net936;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire net935;
 wire _03749_;
 wire net934;
 wire _03751_;
 wire _03752_;
 wire net933;
 wire net932;
 wire net931;
 wire _03756_;
 wire net930;
 wire net929;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire net928;
 wire net927;
 wire _03764_;
 wire _03765_;
 wire net926;
 wire _03767_;
 wire net925;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire net924;
 wire net923;
 wire net922;
 wire _03775_;
 wire net921;
 wire net920;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire net919;
 wire _03783_;
 wire net918;
 wire _03785_;
 wire _03786_;
 wire net917;
 wire net916;
 wire net915;
 wire _03790_;
 wire net914;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire net913;
 wire _03796_;
 wire net912;
 wire _03798_;
 wire _03799_;
 wire net911;
 wire _03801_;
 wire net910;
 wire net909;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire net908;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire net907;
 wire _03812_;
 wire net906;
 wire _03814_;
 wire net905;
 wire _03816_;
 wire _03817_;
 wire net904;
 wire _03819_;
 wire net903;
 wire net902;
 wire net901;
 wire net900;
 wire _03824_;
 wire net899;
 wire _03826_;
 wire net898;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire net897;
 wire net896;
 wire net895;
 wire net894;
 wire _03836_;
 wire _03837_;
 wire net893;
 wire _03839_;
 wire net892;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire net891;
 wire net890;
 wire net889;
 wire _03847_;
 wire net888;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire net887;
 wire net886;
 wire net885;
 wire net884;
 wire _03857_;
 wire net883;
 wire _03859_;
 wire net882;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire net881;
 wire net880;
 wire net879;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire net878;
 wire net877;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire net876;
 wire net875;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire net874;
 wire _03889_;
 wire _03890_;
 wire net873;
 wire net872;
 wire _03893_;
 wire net871;
 wire _03895_;
 wire net870;
 wire _03897_;
 wire net869;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire net868;
 wire _03903_;
 wire net867;
 wire net866;
 wire net865;
 wire net864;
 wire net863;
 wire net862;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire net861;
 wire net860;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire net859;
 wire net858;
 wire net857;
 wire net856;
 wire net855;
 wire net854;
 wire _03924_;
 wire _03925_;
 wire net853;
 wire net852;
 wire net851;
 wire net850;
 wire net849;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire net848;
 wire _03937_;
 wire net847;
 wire net846;
 wire net845;
 wire net844;
 wire net843;
 wire _03943_;
 wire net842;
 wire net841;
 wire net840;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire net839;
 wire _03951_;
 wire _03952_;
 wire net838;
 wire net837;
 wire _03955_;
 wire net836;
 wire net835;
 wire _03958_;
 wire net834;
 wire net833;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire net832;
 wire net831;
 wire net830;
 wire net829;
 wire net828;
 wire _03970_;
 wire net827;
 wire _03972_;
 wire _03973_;
 wire net826;
 wire net825;
 wire net824;
 wire net823;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire net822;
 wire net821;
 wire net820;
 wire net819;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire net818;
 wire net817;
 wire net816;
 wire net815;
 wire net814;
 wire _03995_;
 wire net813;
 wire _03997_;
 wire _03998_;
 wire net812;
 wire _04000_;
 wire net811;
 wire net810;
 wire net809;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire net808;
 wire _04009_;
 wire net807;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire net806;
 wire net805;
 wire net804;
 wire net803;
 wire net802;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire net801;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire net800;
 wire net799;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire net798;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire net797;
 wire _04052_;
 wire _04053_;
 wire net796;
 wire _04055_;
 wire net795;
 wire net794;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire net793;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire net792;
 wire net791;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire net790;
 wire _04103_;
 wire _04104_;
 wire net789;
 wire _04106_;
 wire net788;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire net787;
 wire _04115_;
 wire net786;
 wire net785;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire net784;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire net783;
 wire net782;
 wire net781;
 wire net780;
 wire net779;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire net778;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire net777;
 wire net776;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire net775;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire net774;
 wire _04168_;
 wire _04169_;
 wire net773;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire net772;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire net771;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire net770;
 wire net769;
 wire _04186_;
 wire _04187_;
 wire net768;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire net767;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire net766;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire net765;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire net764;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire net763;
 wire net762;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire net761;
 wire _04235_;
 wire _04236_;
 wire net760;
 wire _04238_;
 wire net759;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire net758;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire net757;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire net756;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire net755;
 wire _04278_;
 wire net754;
 wire _04280_;
 wire _04281_;
 wire net753;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire net752;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire net751;
 wire net750;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire net749;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire net748;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire net747;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire net746;
 wire net745;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire net744;
 wire _04352_;
 wire _04353_;
 wire net743;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire net742;
 wire _04391_;
 wire _04392_;
 wire net741;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire net740;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire net739;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire net738;
 wire _04429_;
 wire net737;
 wire net736;
 wire _04432_;
 wire net735;
 wire _04434_;
 wire net734;
 wire _04436_;
 wire net733;
 wire net732;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire net731;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire net730;
 wire net729;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire net728;
 wire net727;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire net726;
 wire net725;
 wire _04480_;
 wire _04481_;
 wire net724;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire net723;
 wire _04488_;
 wire net722;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire net721;
 wire net720;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire net719;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire net718;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire net717;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire net716;
 wire _04550_;
 wire net715;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire net714;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire net713;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire net712;
 wire _04600_;
 wire net711;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire net710;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire net709;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire net708;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire net707;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire net706;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire net705;
 wire _04736_;
 wire net704;
 wire _04738_;
 wire net703;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire net702;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire net701;
 wire _04780_;
 wire net700;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire net699;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire net698;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire net697;
 wire _04829_;
 wire _04830_;
 wire net696;
 wire _04832_;
 wire net695;
 wire _04834_;
 wire net694;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire net693;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire net692;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire net691;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire net690;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire net689;
 wire _04979_;
 wire _04980_;
 wire net688;
 wire _04982_;
 wire net687;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire net686;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire net685;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire net684;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire net683;
 wire _05036_;
 wire net682;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire net681;
 wire _05063_;
 wire _05064_;
 wire net680;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire net679;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire net678;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire net677;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire net676;
 wire _05120_;
 wire net675;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire net674;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire net673;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire net672;
 wire _05177_;
 wire net671;
 wire _05179_;
 wire _05180_;
 wire net670;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire net669;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire net668;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire net667;
 wire _05205_;
 wire _05206_;
 wire net666;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire net665;
 wire net664;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire net663;
 wire _05225_;
 wire net662;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire net661;
 wire _05236_;
 wire _05237_;
 wire net660;
 wire _05239_;
 wire net659;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire net658;
 wire net657;
 wire _05279_;
 wire _05280_;
 wire net656;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire net655;
 wire _05290_;
 wire _05291_;
 wire net654;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire net653;
 wire net652;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire net651;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire net650;
 wire _05333_;
 wire net649;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire net648;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire net647;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire net646;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire net645;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire net644;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire net643;
 wire net642;
 wire _05423_;
 wire net641;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire net640;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire net639;
 wire _05436_;
 wire _05437_;
 wire net638;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire net637;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire net636;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire net635;
 wire _05455_;
 wire _05456_;
 wire net634;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire net633;
 wire net632;
 wire _05498_;
 wire net631;
 wire _05500_;
 wire net630;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire net629;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire net628;
 wire net627;
 wire _05515_;
 wire _05516_;
 wire net626;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire net625;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire net624;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire net623;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire net622;
 wire _05563_;
 wire net621;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire net620;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire net619;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire net618;
 wire _05582_;
 wire _05583_;
 wire net617;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire net616;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire net615;
 wire _05641_;
 wire net614;
 wire net613;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire net612;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire net611;
 wire _05656_;
 wire net610;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire net609;
 wire _05664_;
 wire _05665_;
 wire net608;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire net607;
 wire _05671_;
 wire net606;
 wire _05673_;
 wire net605;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire net604;
 wire _05680_;
 wire net603;
 wire _05682_;
 wire net602;
 wire _05684_;
 wire net601;
 wire _05686_;
 wire net600;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire net599;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire net598;
 wire net597;
 wire net596;
 wire net595;
 wire net594;
 wire net593;
 wire net592;
 wire net591;
 wire net590;
 wire net589;
 wire _05720_;
 wire net588;
 wire net587;
 wire net586;
 wire _05724_;
 wire net585;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire net584;
 wire net583;
 wire net582;
 wire net581;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire net580;
 wire net579;
 wire net578;
 wire net577;
 wire _05746_;
 wire net576;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire net575;
 wire net574;
 wire net573;
 wire net572;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire net571;
 wire net570;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire net569;
 wire net568;
 wire net567;
 wire _05767_;
 wire _05768_;
 wire net566;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire net565;
 wire _05776_;
 wire net564;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire net563;
 wire net562;
 wire _05788_;
 wire net561;
 wire _05790_;
 wire _05791_;
 wire net560;
 wire _05793_;
 wire net559;
 wire _05795_;
 wire net558;
 wire net557;
 wire _05798_;
 wire net556;
 wire _05800_;
 wire net555;
 wire net554;
 wire _05803_;
 wire _05804_;
 wire net553;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire net552;
 wire net550;
 wire net551;
 wire _05814_;
 wire net549;
 wire net548;
 wire net547;
 wire _05818_;
 wire net546;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire net545;
 wire net544;
 wire net543;
 wire net542;
 wire _05828_;
 wire _05829_;
 wire net541;
 wire net540;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire net539;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire net538;
 wire _05842_;
 wire net537;
 wire _05844_;
 wire net536;
 wire net535;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire net534;
 wire _05852_;
 wire _05853_;
 wire net533;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire net532;
 wire _05870_;
 wire _05871_;
 wire net531;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire net530;
 wire _05878_;
 wire _05879_;
 wire net529;
 wire net528;
 wire net527;
 wire _05883_;
 wire _05884_;
 wire net526;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire net525;
 wire _05890_;
 wire _05891_;
 wire net524;
 wire net523;
 wire _05894_;
 wire net522;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire net521;
 wire net520;
 wire net519;
 wire _05902_;
 wire net518;
 wire net517;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire net516;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire net515;
 wire _05914_;
 wire net514;
 wire net513;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire net512;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire net511;
 wire _05942_;
 wire net510;
 wire _05944_;
 wire net509;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire net508;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire net507;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire net506;
 wire net505;
 wire net504;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire net503;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire net502;
 wire _06001_;
 wire net501;
 wire _06003_;
 wire _06004_;
 wire net500;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire net499;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire net498;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire net497;
 wire _06022_;
 wire net496;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire net495;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire net494;
 wire net493;
 wire net492;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire net491;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire net490;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire net489;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire net488;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire net487;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire net486;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire net485;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire net484;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire net483;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire net482;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire net481;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire net480;
 wire _06191_;
 wire net479;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire net478;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire net477;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire net476;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire net475;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire net474;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire net473;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire net472;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire net471;
 wire _06607_;
 wire net470;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire net469;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire net468;
 wire _06780_;
 wire net467;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire net466;
 wire _06788_;
 wire _06789_;
 wire net465;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire net464;
 wire _06796_;
 wire _06797_;
 wire net463;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire net462;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire net461;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire net460;
 wire _06843_;
 wire _06844_;
 wire net459;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire net458;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire net457;
 wire net456;
 wire net455;
 wire net454;
 wire net453;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire net452;
 wire net451;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire net450;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire net449;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire net448;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire net447;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire net446;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire net445;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire net444;
 wire _07066_;
 wire net443;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire net442;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire net441;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire net440;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire net439;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire net438;
 wire _07112_;
 wire net437;
 wire _07114_;
 wire net436;
 wire _07116_;
 wire _07117_;
 wire net435;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire net434;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire net433;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire net432;
 wire _07178_;
 wire _07179_;
 wire net431;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire net430;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire net429;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire net428;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire net427;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire net426;
 wire _07232_;
 wire _07233_;
 wire net425;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire net424;
 wire _07240_;
 wire net423;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire net422;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire net421;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire net420;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire net419;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire net418;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire net417;
 wire _07315_;
 wire _07316_;
 wire net416;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire net415;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire net414;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire net413;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire net412;
 wire net411;
 wire _07393_;
 wire net410;
 wire _07395_;
 wire _07396_;
 wire net409;
 wire _07398_;
 wire net408;
 wire net407;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire net406;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire net405;
 wire net404;
 wire _07414_;
 wire net403;
 wire net402;
 wire net401;
 wire net400;
 wire net399;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire net398;
 wire _07426_;
 wire _07427_;
 wire net397;
 wire net396;
 wire _07430_;
 wire _07431_;
 wire net395;
 wire net394;
 wire _07434_;
 wire net393;
 wire net392;
 wire net391;
 wire _07438_;
 wire net390;
 wire net389;
 wire _07441_;
 wire _07442_;
 wire net388;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire net387;
 wire net386;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire net385;
 wire net384;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire net383;
 wire net382;
 wire _07465_;
 wire net381;
 wire _07467_;
 wire _07468_;
 wire net380;
 wire net379;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire net378;
 wire net377;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire net376;
 wire net375;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire net374;
 wire _07491_;
 wire _07492_;
 wire net373;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire net372;
 wire net371;
 wire _07501_;
 wire _07502_;
 wire net370;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire net369;
 wire net368;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire net367;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire net366;
 wire net365;
 wire net364;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire net363;
 wire net362;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire net361;
 wire net360;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire net359;
 wire net358;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire net357;
 wire net356;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire net355;
 wire net354;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire net353;
 wire net352;
 wire net351;
 wire _07568_;
 wire _07569_;
 wire net350;
 wire net349;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire net348;
 wire net347;
 wire _07579_;
 wire net346;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire net345;
 wire net344;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire net343;
 wire net342;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire net341;
 wire net340;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire net339;
 wire net338;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire net337;
 wire net336;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire net335;
 wire net334;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire net333;
 wire net332;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire net331;
 wire net330;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire net329;
 wire net328;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire net327;
 wire net326;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire net325;
 wire net324;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire net323;
 wire net322;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire net321;
 wire net320;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire net319;
 wire net318;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire net317;
 wire net316;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire net315;
 wire _07748_;
 wire net314;
 wire net313;
 wire net312;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire net311;
 wire _07761_;
 wire _07762_;
 wire net310;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire net309;
 wire _07773_;
 wire _07774_;
 wire net308;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire net307;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire net306;
 wire _07789_;
 wire _07790_;
 wire net305;
 wire _07792_;
 wire net304;
 wire _07794_;
 wire _07795_;
 wire net303;
 wire _07797_;
 wire net302;
 wire net301;
 wire net300;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire net299;
 wire _07805_;
 wire _07806_;
 wire net298;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire net297;
 wire _07814_;
 wire net296;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire net295;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire net294;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire net293;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire net292;
 wire _07838_;
 wire net291;
 wire _07840_;
 wire _07841_;
 wire net290;
 wire _07843_;
 wire net289;
 wire net288;
 wire net287;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire net286;
 wire _07856_;
 wire _07857_;
 wire net285;
 wire _07859_;
 wire _07860_;
 wire net284;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire net283;
 wire _07869_;
 wire _07870_;
 wire net282;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire net281;
 wire net280;
 wire net279;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire net278;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire net277;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire net276;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire net275;
 wire _07906_;
 wire net274;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire net273;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire net272;
 wire _07926_;
 wire net271;
 wire net270;
 wire _07929_;
 wire _07930_;
 wire net269;
 wire _07932_;
 wire net268;
 wire net267;
 wire net266;
 wire net265;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire net264;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire net263;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire net262;
 wire net261;
 wire net260;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire net259;
 wire _07981_;
 wire _07982_;
 wire net258;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire net257;
 wire _07993_;
 wire _07994_;
 wire net256;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire net255;
 wire net254;
 wire net253;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire net252;
 wire _08015_;
 wire _08016_;
 wire net251;
 wire _08018_;
 wire net250;
 wire _08020_;
 wire net249;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire net248;
 wire _08028_;
 wire _08029_;
 wire net247;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire net246;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire net245;
 wire net244;
 wire net243;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire net242;
 wire net241;
 wire net240;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire net239;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire net238;
 wire net237;
 wire _08094_;
 wire _08095_;
 wire net236;
 wire net235;
 wire net234;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire net233;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire net232;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire net231;
 wire net230;
 wire net229;
 wire _08134_;
 wire net228;
 wire _08136_;
 wire net227;
 wire _08138_;
 wire net226;
 wire _08140_;
 wire net225;
 wire _08142_;
 wire net224;
 wire _08144_;
 wire net223;
 wire _08146_;
 wire net222;
 wire _08148_;
 wire net221;
 wire net220;
 wire _08151_;
 wire net219;
 wire _08153_;
 wire net218;
 wire net217;
 wire _08156_;
 wire net216;
 wire _08158_;
 wire _08159_;
 wire net215;
 wire _08161_;
 wire net214;
 wire _08163_;
 wire _08164_;
 wire net213;
 wire _08166_;
 wire net212;
 wire _08168_;
 wire net211;
 wire _08170_;
 wire net210;
 wire _08172_;
 wire net209;
 wire _08174_;
 wire net208;
 wire _08176_;
 wire net207;
 wire _08178_;
 wire net206;
 wire _08180_;
 wire net205;
 wire _08182_;
 wire net204;
 wire _08184_;
 wire net203;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire net202;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire net201;
 wire net200;
 wire net199;
 wire _08196_;
 wire _08197_;
 wire net198;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire net197;
 wire _08203_;
 wire net196;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire net195;
 wire _08212_;
 wire _08213_;
 wire net194;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire net193;
 wire net192;
 wire net191;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire net190;
 wire _08246_;
 wire _08247_;
 wire net189;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire net188;
 wire _08258_;
 wire _08259_;
 wire net187;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire net186;
 wire net185;
 wire net184;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire net183;
 wire _08284_;
 wire _08285_;
 wire net182;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire net181;
 wire _08296_;
 wire _08297_;
 wire net180;
 wire net179;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire net178;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire net177;
 wire net176;
 wire net175;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire net174;
 wire _08325_;
 wire _08326_;
 wire net173;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire net172;
 wire _08337_;
 wire _08338_;
 wire net171;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire net140;
 wire net139;
 wire net138;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire net137;
 wire _08363_;
 wire _08364_;
 wire net136;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire net135;
 wire _08375_;
 wire _08376_;
 wire net134;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire net133;
 wire _08389_;
 wire net132;
 wire net131;
 wire net130;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire net129;
 wire _08402_;
 wire _08403_;
 wire net128;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire net127;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire net126;
 wire _08415_;
 wire _08416_;
 wire net125;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire net124;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire net123;
 wire net122;
 wire net121;
 wire _08433_;
 wire _08434_;
 wire net120;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire net119;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire net118;
 wire _08447_;
 wire _08448_;
 wire net117;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire net116;
 wire _08470_;
 wire net115;
 wire net114;
 wire _08473_;
 wire _08474_;
 wire net113;
 wire net112;
 wire net111;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire net110;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire net109;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire net108;
 wire _08511_;
 wire _08512_;
 wire net107;
 wire net106;
 wire net105;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire \dp.ISRmux.d0[10] ;
 wire \dp.ISRmux.d0[11] ;
 wire \dp.ISRmux.d0[12] ;
 wire \dp.ISRmux.d0[13] ;
 wire \dp.ISRmux.d0[14] ;
 wire \dp.ISRmux.d0[15] ;
 wire \dp.ISRmux.d0[16] ;
 wire \dp.ISRmux.d0[17] ;
 wire \dp.ISRmux.d0[18] ;
 wire \dp.ISRmux.d0[19] ;
 wire \dp.ISRmux.d0[20] ;
 wire \dp.ISRmux.d0[21] ;
 wire \dp.ISRmux.d0[22] ;
 wire \dp.ISRmux.d0[23] ;
 wire \dp.ISRmux.d0[24] ;
 wire \dp.ISRmux.d0[25] ;
 wire \dp.ISRmux.d0[26] ;
 wire \dp.ISRmux.d0[27] ;
 wire \dp.ISRmux.d0[28] ;
 wire \dp.ISRmux.d0[29] ;
 wire \dp.ISRmux.d0[2] ;
 wire \dp.ISRmux.d0[30] ;
 wire \dp.ISRmux.d0[31] ;
 wire \dp.ISRmux.d0[3] ;
 wire \dp.ISRmux.d0[4] ;
 wire \dp.ISRmux.d0[5] ;
 wire \dp.ISRmux.d0[6] ;
 wire \dp.ISRmux.d0[7] ;
 wire \dp.ISRmux.d0[8] ;
 wire \dp.ISRmux.d0[9] ;
 wire \dp.rf.rf[0][0] ;
 wire \dp.rf.rf[0][10] ;
 wire \dp.rf.rf[0][11] ;
 wire \dp.rf.rf[0][12] ;
 wire \dp.rf.rf[0][13] ;
 wire \dp.rf.rf[0][14] ;
 wire \dp.rf.rf[0][15] ;
 wire \dp.rf.rf[0][16] ;
 wire \dp.rf.rf[0][18] ;
 wire \dp.rf.rf[0][1] ;
 wire \dp.rf.rf[0][20] ;
 wire \dp.rf.rf[0][21] ;
 wire \dp.rf.rf[0][22] ;
 wire \dp.rf.rf[0][23] ;
 wire \dp.rf.rf[0][24] ;
 wire \dp.rf.rf[0][25] ;
 wire \dp.rf.rf[0][26] ;
 wire \dp.rf.rf[0][27] ;
 wire \dp.rf.rf[0][28] ;
 wire \dp.rf.rf[0][29] ;
 wire \dp.rf.rf[0][2] ;
 wire \dp.rf.rf[0][30] ;
 wire \dp.rf.rf[0][31] ;
 wire \dp.rf.rf[0][3] ;
 wire \dp.rf.rf[0][4] ;
 wire \dp.rf.rf[0][5] ;
 wire \dp.rf.rf[0][6] ;
 wire \dp.rf.rf[0][7] ;
 wire \dp.rf.rf[0][8] ;
 wire \dp.rf.rf[0][9] ;
 wire \dp.rf.rf[10][0] ;
 wire \dp.rf.rf[10][10] ;
 wire \dp.rf.rf[10][11] ;
 wire \dp.rf.rf[10][12] ;
 wire \dp.rf.rf[10][13] ;
 wire \dp.rf.rf[10][14] ;
 wire \dp.rf.rf[10][15] ;
 wire \dp.rf.rf[10][16] ;
 wire \dp.rf.rf[10][17] ;
 wire \dp.rf.rf[10][18] ;
 wire \dp.rf.rf[10][19] ;
 wire \dp.rf.rf[10][1] ;
 wire \dp.rf.rf[10][20] ;
 wire \dp.rf.rf[10][21] ;
 wire \dp.rf.rf[10][22] ;
 wire \dp.rf.rf[10][23] ;
 wire \dp.rf.rf[10][24] ;
 wire \dp.rf.rf[10][25] ;
 wire \dp.rf.rf[10][26] ;
 wire \dp.rf.rf[10][27] ;
 wire \dp.rf.rf[10][28] ;
 wire \dp.rf.rf[10][29] ;
 wire \dp.rf.rf[10][2] ;
 wire \dp.rf.rf[10][30] ;
 wire \dp.rf.rf[10][31] ;
 wire \dp.rf.rf[10][3] ;
 wire \dp.rf.rf[10][4] ;
 wire \dp.rf.rf[10][5] ;
 wire \dp.rf.rf[10][6] ;
 wire \dp.rf.rf[10][7] ;
 wire \dp.rf.rf[10][8] ;
 wire \dp.rf.rf[10][9] ;
 wire \dp.rf.rf[11][0] ;
 wire \dp.rf.rf[11][10] ;
 wire \dp.rf.rf[11][11] ;
 wire \dp.rf.rf[11][12] ;
 wire \dp.rf.rf[11][13] ;
 wire \dp.rf.rf[11][14] ;
 wire \dp.rf.rf[11][15] ;
 wire \dp.rf.rf[11][16] ;
 wire \dp.rf.rf[11][17] ;
 wire \dp.rf.rf[11][18] ;
 wire \dp.rf.rf[11][19] ;
 wire \dp.rf.rf[11][1] ;
 wire \dp.rf.rf[11][20] ;
 wire \dp.rf.rf[11][21] ;
 wire \dp.rf.rf[11][22] ;
 wire \dp.rf.rf[11][23] ;
 wire \dp.rf.rf[11][24] ;
 wire \dp.rf.rf[11][25] ;
 wire \dp.rf.rf[11][26] ;
 wire \dp.rf.rf[11][27] ;
 wire \dp.rf.rf[11][28] ;
 wire \dp.rf.rf[11][29] ;
 wire \dp.rf.rf[11][2] ;
 wire \dp.rf.rf[11][30] ;
 wire \dp.rf.rf[11][31] ;
 wire \dp.rf.rf[11][3] ;
 wire \dp.rf.rf[11][4] ;
 wire \dp.rf.rf[11][5] ;
 wire \dp.rf.rf[11][6] ;
 wire \dp.rf.rf[11][7] ;
 wire \dp.rf.rf[11][8] ;
 wire \dp.rf.rf[11][9] ;
 wire \dp.rf.rf[12][0] ;
 wire \dp.rf.rf[12][10] ;
 wire \dp.rf.rf[12][11] ;
 wire \dp.rf.rf[12][12] ;
 wire \dp.rf.rf[12][13] ;
 wire \dp.rf.rf[12][14] ;
 wire \dp.rf.rf[12][15] ;
 wire \dp.rf.rf[12][16] ;
 wire \dp.rf.rf[12][17] ;
 wire \dp.rf.rf[12][18] ;
 wire \dp.rf.rf[12][19] ;
 wire \dp.rf.rf[12][1] ;
 wire \dp.rf.rf[12][20] ;
 wire \dp.rf.rf[12][21] ;
 wire \dp.rf.rf[12][22] ;
 wire \dp.rf.rf[12][23] ;
 wire \dp.rf.rf[12][24] ;
 wire \dp.rf.rf[12][25] ;
 wire \dp.rf.rf[12][26] ;
 wire \dp.rf.rf[12][27] ;
 wire \dp.rf.rf[12][28] ;
 wire \dp.rf.rf[12][29] ;
 wire \dp.rf.rf[12][2] ;
 wire \dp.rf.rf[12][30] ;
 wire \dp.rf.rf[12][31] ;
 wire \dp.rf.rf[12][3] ;
 wire \dp.rf.rf[12][4] ;
 wire \dp.rf.rf[12][5] ;
 wire \dp.rf.rf[12][6] ;
 wire \dp.rf.rf[12][7] ;
 wire \dp.rf.rf[12][8] ;
 wire \dp.rf.rf[12][9] ;
 wire \dp.rf.rf[13][0] ;
 wire \dp.rf.rf[13][10] ;
 wire \dp.rf.rf[13][11] ;
 wire \dp.rf.rf[13][12] ;
 wire \dp.rf.rf[13][13] ;
 wire \dp.rf.rf[13][14] ;
 wire \dp.rf.rf[13][15] ;
 wire \dp.rf.rf[13][16] ;
 wire \dp.rf.rf[13][17] ;
 wire \dp.rf.rf[13][18] ;
 wire \dp.rf.rf[13][19] ;
 wire \dp.rf.rf[13][1] ;
 wire \dp.rf.rf[13][20] ;
 wire \dp.rf.rf[13][21] ;
 wire \dp.rf.rf[13][22] ;
 wire \dp.rf.rf[13][23] ;
 wire \dp.rf.rf[13][24] ;
 wire \dp.rf.rf[13][25] ;
 wire \dp.rf.rf[13][26] ;
 wire \dp.rf.rf[13][27] ;
 wire \dp.rf.rf[13][28] ;
 wire \dp.rf.rf[13][29] ;
 wire \dp.rf.rf[13][2] ;
 wire \dp.rf.rf[13][30] ;
 wire \dp.rf.rf[13][31] ;
 wire \dp.rf.rf[13][3] ;
 wire \dp.rf.rf[13][4] ;
 wire \dp.rf.rf[13][5] ;
 wire \dp.rf.rf[13][6] ;
 wire \dp.rf.rf[13][7] ;
 wire \dp.rf.rf[13][8] ;
 wire \dp.rf.rf[13][9] ;
 wire \dp.rf.rf[14][0] ;
 wire \dp.rf.rf[14][10] ;
 wire \dp.rf.rf[14][11] ;
 wire \dp.rf.rf[14][12] ;
 wire \dp.rf.rf[14][13] ;
 wire \dp.rf.rf[14][14] ;
 wire \dp.rf.rf[14][15] ;
 wire \dp.rf.rf[14][16] ;
 wire \dp.rf.rf[14][17] ;
 wire \dp.rf.rf[14][18] ;
 wire \dp.rf.rf[14][19] ;
 wire \dp.rf.rf[14][1] ;
 wire \dp.rf.rf[14][20] ;
 wire \dp.rf.rf[14][21] ;
 wire \dp.rf.rf[14][22] ;
 wire \dp.rf.rf[14][23] ;
 wire \dp.rf.rf[14][24] ;
 wire \dp.rf.rf[14][25] ;
 wire \dp.rf.rf[14][26] ;
 wire \dp.rf.rf[14][27] ;
 wire \dp.rf.rf[14][28] ;
 wire \dp.rf.rf[14][29] ;
 wire \dp.rf.rf[14][2] ;
 wire \dp.rf.rf[14][30] ;
 wire \dp.rf.rf[14][31] ;
 wire \dp.rf.rf[14][3] ;
 wire \dp.rf.rf[14][4] ;
 wire \dp.rf.rf[14][5] ;
 wire \dp.rf.rf[14][6] ;
 wire \dp.rf.rf[14][7] ;
 wire \dp.rf.rf[14][8] ;
 wire \dp.rf.rf[14][9] ;
 wire \dp.rf.rf[15][0] ;
 wire \dp.rf.rf[15][10] ;
 wire \dp.rf.rf[15][11] ;
 wire \dp.rf.rf[15][12] ;
 wire \dp.rf.rf[15][13] ;
 wire \dp.rf.rf[15][14] ;
 wire \dp.rf.rf[15][15] ;
 wire \dp.rf.rf[15][16] ;
 wire \dp.rf.rf[15][17] ;
 wire \dp.rf.rf[15][18] ;
 wire \dp.rf.rf[15][19] ;
 wire \dp.rf.rf[15][1] ;
 wire \dp.rf.rf[15][20] ;
 wire \dp.rf.rf[15][21] ;
 wire \dp.rf.rf[15][22] ;
 wire \dp.rf.rf[15][23] ;
 wire \dp.rf.rf[15][24] ;
 wire \dp.rf.rf[15][25] ;
 wire \dp.rf.rf[15][26] ;
 wire \dp.rf.rf[15][27] ;
 wire \dp.rf.rf[15][28] ;
 wire \dp.rf.rf[15][29] ;
 wire \dp.rf.rf[15][2] ;
 wire \dp.rf.rf[15][30] ;
 wire \dp.rf.rf[15][31] ;
 wire \dp.rf.rf[15][3] ;
 wire \dp.rf.rf[15][4] ;
 wire \dp.rf.rf[15][5] ;
 wire \dp.rf.rf[15][6] ;
 wire \dp.rf.rf[15][7] ;
 wire \dp.rf.rf[15][8] ;
 wire \dp.rf.rf[15][9] ;
 wire \dp.rf.rf[16][0] ;
 wire \dp.rf.rf[16][10] ;
 wire \dp.rf.rf[16][11] ;
 wire \dp.rf.rf[16][12] ;
 wire \dp.rf.rf[16][13] ;
 wire \dp.rf.rf[16][14] ;
 wire \dp.rf.rf[16][15] ;
 wire \dp.rf.rf[16][16] ;
 wire \dp.rf.rf[16][17] ;
 wire \dp.rf.rf[16][18] ;
 wire \dp.rf.rf[16][19] ;
 wire \dp.rf.rf[16][1] ;
 wire \dp.rf.rf[16][20] ;
 wire \dp.rf.rf[16][21] ;
 wire \dp.rf.rf[16][22] ;
 wire \dp.rf.rf[16][23] ;
 wire \dp.rf.rf[16][24] ;
 wire \dp.rf.rf[16][25] ;
 wire \dp.rf.rf[16][26] ;
 wire \dp.rf.rf[16][27] ;
 wire \dp.rf.rf[16][28] ;
 wire \dp.rf.rf[16][29] ;
 wire \dp.rf.rf[16][2] ;
 wire \dp.rf.rf[16][30] ;
 wire \dp.rf.rf[16][31] ;
 wire \dp.rf.rf[16][3] ;
 wire \dp.rf.rf[16][4] ;
 wire \dp.rf.rf[16][5] ;
 wire \dp.rf.rf[16][6] ;
 wire \dp.rf.rf[16][7] ;
 wire \dp.rf.rf[16][8] ;
 wire \dp.rf.rf[16][9] ;
 wire \dp.rf.rf[17][0] ;
 wire \dp.rf.rf[17][10] ;
 wire \dp.rf.rf[17][11] ;
 wire \dp.rf.rf[17][12] ;
 wire \dp.rf.rf[17][13] ;
 wire \dp.rf.rf[17][14] ;
 wire \dp.rf.rf[17][15] ;
 wire \dp.rf.rf[17][16] ;
 wire \dp.rf.rf[17][17] ;
 wire \dp.rf.rf[17][18] ;
 wire \dp.rf.rf[17][19] ;
 wire \dp.rf.rf[17][1] ;
 wire \dp.rf.rf[17][20] ;
 wire \dp.rf.rf[17][21] ;
 wire \dp.rf.rf[17][22] ;
 wire \dp.rf.rf[17][23] ;
 wire \dp.rf.rf[17][24] ;
 wire \dp.rf.rf[17][25] ;
 wire \dp.rf.rf[17][26] ;
 wire \dp.rf.rf[17][27] ;
 wire \dp.rf.rf[17][28] ;
 wire \dp.rf.rf[17][29] ;
 wire \dp.rf.rf[17][2] ;
 wire \dp.rf.rf[17][30] ;
 wire \dp.rf.rf[17][31] ;
 wire \dp.rf.rf[17][3] ;
 wire \dp.rf.rf[17][4] ;
 wire \dp.rf.rf[17][5] ;
 wire \dp.rf.rf[17][6] ;
 wire \dp.rf.rf[17][7] ;
 wire \dp.rf.rf[17][8] ;
 wire \dp.rf.rf[17][9] ;
 wire \dp.rf.rf[18][0] ;
 wire \dp.rf.rf[18][10] ;
 wire \dp.rf.rf[18][11] ;
 wire \dp.rf.rf[18][12] ;
 wire \dp.rf.rf[18][13] ;
 wire \dp.rf.rf[18][14] ;
 wire \dp.rf.rf[18][15] ;
 wire \dp.rf.rf[18][16] ;
 wire \dp.rf.rf[18][17] ;
 wire \dp.rf.rf[18][18] ;
 wire \dp.rf.rf[18][19] ;
 wire \dp.rf.rf[18][1] ;
 wire \dp.rf.rf[18][20] ;
 wire \dp.rf.rf[18][21] ;
 wire \dp.rf.rf[18][22] ;
 wire \dp.rf.rf[18][23] ;
 wire \dp.rf.rf[18][24] ;
 wire \dp.rf.rf[18][25] ;
 wire \dp.rf.rf[18][26] ;
 wire \dp.rf.rf[18][27] ;
 wire \dp.rf.rf[18][28] ;
 wire \dp.rf.rf[18][29] ;
 wire \dp.rf.rf[18][2] ;
 wire \dp.rf.rf[18][30] ;
 wire \dp.rf.rf[18][31] ;
 wire \dp.rf.rf[18][3] ;
 wire \dp.rf.rf[18][4] ;
 wire \dp.rf.rf[18][5] ;
 wire \dp.rf.rf[18][6] ;
 wire \dp.rf.rf[18][7] ;
 wire \dp.rf.rf[18][8] ;
 wire \dp.rf.rf[18][9] ;
 wire \dp.rf.rf[19][0] ;
 wire \dp.rf.rf[19][10] ;
 wire \dp.rf.rf[19][11] ;
 wire \dp.rf.rf[19][12] ;
 wire \dp.rf.rf[19][13] ;
 wire \dp.rf.rf[19][14] ;
 wire \dp.rf.rf[19][15] ;
 wire \dp.rf.rf[19][16] ;
 wire \dp.rf.rf[19][17] ;
 wire \dp.rf.rf[19][18] ;
 wire \dp.rf.rf[19][19] ;
 wire \dp.rf.rf[19][1] ;
 wire \dp.rf.rf[19][20] ;
 wire \dp.rf.rf[19][21] ;
 wire \dp.rf.rf[19][22] ;
 wire \dp.rf.rf[19][23] ;
 wire \dp.rf.rf[19][24] ;
 wire \dp.rf.rf[19][25] ;
 wire \dp.rf.rf[19][26] ;
 wire \dp.rf.rf[19][27] ;
 wire \dp.rf.rf[19][28] ;
 wire \dp.rf.rf[19][29] ;
 wire \dp.rf.rf[19][2] ;
 wire \dp.rf.rf[19][30] ;
 wire \dp.rf.rf[19][31] ;
 wire \dp.rf.rf[19][3] ;
 wire \dp.rf.rf[19][4] ;
 wire \dp.rf.rf[19][5] ;
 wire \dp.rf.rf[19][6] ;
 wire \dp.rf.rf[19][7] ;
 wire \dp.rf.rf[19][8] ;
 wire \dp.rf.rf[19][9] ;
 wire \dp.rf.rf[1][0] ;
 wire \dp.rf.rf[1][10] ;
 wire \dp.rf.rf[1][11] ;
 wire \dp.rf.rf[1][12] ;
 wire \dp.rf.rf[1][13] ;
 wire \dp.rf.rf[1][14] ;
 wire \dp.rf.rf[1][15] ;
 wire \dp.rf.rf[1][16] ;
 wire \dp.rf.rf[1][17] ;
 wire \dp.rf.rf[1][18] ;
 wire \dp.rf.rf[1][19] ;
 wire \dp.rf.rf[1][1] ;
 wire \dp.rf.rf[1][20] ;
 wire \dp.rf.rf[1][21] ;
 wire \dp.rf.rf[1][22] ;
 wire \dp.rf.rf[1][23] ;
 wire \dp.rf.rf[1][24] ;
 wire \dp.rf.rf[1][25] ;
 wire \dp.rf.rf[1][26] ;
 wire \dp.rf.rf[1][27] ;
 wire \dp.rf.rf[1][28] ;
 wire \dp.rf.rf[1][29] ;
 wire \dp.rf.rf[1][2] ;
 wire \dp.rf.rf[1][30] ;
 wire \dp.rf.rf[1][31] ;
 wire \dp.rf.rf[1][3] ;
 wire \dp.rf.rf[1][4] ;
 wire \dp.rf.rf[1][5] ;
 wire \dp.rf.rf[1][6] ;
 wire \dp.rf.rf[1][7] ;
 wire \dp.rf.rf[1][8] ;
 wire \dp.rf.rf[1][9] ;
 wire \dp.rf.rf[20][0] ;
 wire \dp.rf.rf[20][10] ;
 wire \dp.rf.rf[20][11] ;
 wire \dp.rf.rf[20][12] ;
 wire \dp.rf.rf[20][13] ;
 wire \dp.rf.rf[20][14] ;
 wire \dp.rf.rf[20][15] ;
 wire \dp.rf.rf[20][16] ;
 wire \dp.rf.rf[20][17] ;
 wire \dp.rf.rf[20][18] ;
 wire \dp.rf.rf[20][19] ;
 wire \dp.rf.rf[20][1] ;
 wire \dp.rf.rf[20][20] ;
 wire \dp.rf.rf[20][21] ;
 wire \dp.rf.rf[20][22] ;
 wire \dp.rf.rf[20][23] ;
 wire \dp.rf.rf[20][24] ;
 wire \dp.rf.rf[20][25] ;
 wire \dp.rf.rf[20][26] ;
 wire \dp.rf.rf[20][27] ;
 wire \dp.rf.rf[20][28] ;
 wire \dp.rf.rf[20][29] ;
 wire \dp.rf.rf[20][2] ;
 wire \dp.rf.rf[20][30] ;
 wire \dp.rf.rf[20][31] ;
 wire \dp.rf.rf[20][3] ;
 wire \dp.rf.rf[20][4] ;
 wire \dp.rf.rf[20][5] ;
 wire \dp.rf.rf[20][6] ;
 wire \dp.rf.rf[20][7] ;
 wire \dp.rf.rf[20][8] ;
 wire \dp.rf.rf[20][9] ;
 wire \dp.rf.rf[21][0] ;
 wire \dp.rf.rf[21][10] ;
 wire \dp.rf.rf[21][11] ;
 wire \dp.rf.rf[21][12] ;
 wire \dp.rf.rf[21][13] ;
 wire \dp.rf.rf[21][14] ;
 wire \dp.rf.rf[21][15] ;
 wire \dp.rf.rf[21][16] ;
 wire \dp.rf.rf[21][17] ;
 wire \dp.rf.rf[21][18] ;
 wire \dp.rf.rf[21][19] ;
 wire \dp.rf.rf[21][1] ;
 wire \dp.rf.rf[21][20] ;
 wire \dp.rf.rf[21][21] ;
 wire \dp.rf.rf[21][22] ;
 wire \dp.rf.rf[21][23] ;
 wire \dp.rf.rf[21][24] ;
 wire \dp.rf.rf[21][25] ;
 wire \dp.rf.rf[21][26] ;
 wire \dp.rf.rf[21][27] ;
 wire \dp.rf.rf[21][28] ;
 wire \dp.rf.rf[21][29] ;
 wire \dp.rf.rf[21][2] ;
 wire \dp.rf.rf[21][30] ;
 wire \dp.rf.rf[21][31] ;
 wire \dp.rf.rf[21][3] ;
 wire \dp.rf.rf[21][4] ;
 wire \dp.rf.rf[21][5] ;
 wire \dp.rf.rf[21][6] ;
 wire \dp.rf.rf[21][7] ;
 wire \dp.rf.rf[21][8] ;
 wire \dp.rf.rf[21][9] ;
 wire \dp.rf.rf[22][0] ;
 wire \dp.rf.rf[22][10] ;
 wire \dp.rf.rf[22][11] ;
 wire \dp.rf.rf[22][12] ;
 wire \dp.rf.rf[22][13] ;
 wire \dp.rf.rf[22][14] ;
 wire \dp.rf.rf[22][15] ;
 wire \dp.rf.rf[22][16] ;
 wire \dp.rf.rf[22][17] ;
 wire \dp.rf.rf[22][18] ;
 wire \dp.rf.rf[22][19] ;
 wire \dp.rf.rf[22][1] ;
 wire \dp.rf.rf[22][20] ;
 wire \dp.rf.rf[22][21] ;
 wire \dp.rf.rf[22][22] ;
 wire \dp.rf.rf[22][23] ;
 wire \dp.rf.rf[22][24] ;
 wire \dp.rf.rf[22][25] ;
 wire \dp.rf.rf[22][26] ;
 wire \dp.rf.rf[22][27] ;
 wire \dp.rf.rf[22][28] ;
 wire \dp.rf.rf[22][29] ;
 wire \dp.rf.rf[22][2] ;
 wire \dp.rf.rf[22][30] ;
 wire \dp.rf.rf[22][31] ;
 wire \dp.rf.rf[22][3] ;
 wire \dp.rf.rf[22][4] ;
 wire \dp.rf.rf[22][5] ;
 wire \dp.rf.rf[22][6] ;
 wire \dp.rf.rf[22][7] ;
 wire \dp.rf.rf[22][8] ;
 wire \dp.rf.rf[22][9] ;
 wire \dp.rf.rf[23][0] ;
 wire \dp.rf.rf[23][10] ;
 wire \dp.rf.rf[23][11] ;
 wire \dp.rf.rf[23][12] ;
 wire \dp.rf.rf[23][13] ;
 wire \dp.rf.rf[23][14] ;
 wire \dp.rf.rf[23][15] ;
 wire \dp.rf.rf[23][16] ;
 wire \dp.rf.rf[23][17] ;
 wire \dp.rf.rf[23][18] ;
 wire \dp.rf.rf[23][19] ;
 wire \dp.rf.rf[23][1] ;
 wire \dp.rf.rf[23][20] ;
 wire \dp.rf.rf[23][21] ;
 wire \dp.rf.rf[23][22] ;
 wire \dp.rf.rf[23][23] ;
 wire \dp.rf.rf[23][24] ;
 wire \dp.rf.rf[23][25] ;
 wire \dp.rf.rf[23][26] ;
 wire \dp.rf.rf[23][27] ;
 wire \dp.rf.rf[23][28] ;
 wire \dp.rf.rf[23][29] ;
 wire \dp.rf.rf[23][2] ;
 wire \dp.rf.rf[23][30] ;
 wire \dp.rf.rf[23][31] ;
 wire \dp.rf.rf[23][3] ;
 wire \dp.rf.rf[23][4] ;
 wire \dp.rf.rf[23][5] ;
 wire \dp.rf.rf[23][6] ;
 wire \dp.rf.rf[23][7] ;
 wire \dp.rf.rf[23][8] ;
 wire \dp.rf.rf[23][9] ;
 wire \dp.rf.rf[24][0] ;
 wire \dp.rf.rf[24][10] ;
 wire \dp.rf.rf[24][11] ;
 wire \dp.rf.rf[24][12] ;
 wire \dp.rf.rf[24][13] ;
 wire \dp.rf.rf[24][14] ;
 wire \dp.rf.rf[24][15] ;
 wire \dp.rf.rf[24][16] ;
 wire \dp.rf.rf[24][17] ;
 wire \dp.rf.rf[24][18] ;
 wire \dp.rf.rf[24][19] ;
 wire \dp.rf.rf[24][1] ;
 wire \dp.rf.rf[24][20] ;
 wire \dp.rf.rf[24][21] ;
 wire \dp.rf.rf[24][22] ;
 wire \dp.rf.rf[24][23] ;
 wire \dp.rf.rf[24][24] ;
 wire \dp.rf.rf[24][25] ;
 wire \dp.rf.rf[24][26] ;
 wire \dp.rf.rf[24][27] ;
 wire \dp.rf.rf[24][28] ;
 wire \dp.rf.rf[24][29] ;
 wire \dp.rf.rf[24][2] ;
 wire \dp.rf.rf[24][30] ;
 wire \dp.rf.rf[24][31] ;
 wire \dp.rf.rf[24][3] ;
 wire \dp.rf.rf[24][4] ;
 wire \dp.rf.rf[24][5] ;
 wire \dp.rf.rf[24][6] ;
 wire \dp.rf.rf[24][7] ;
 wire \dp.rf.rf[24][8] ;
 wire \dp.rf.rf[24][9] ;
 wire \dp.rf.rf[25][0] ;
 wire \dp.rf.rf[25][10] ;
 wire \dp.rf.rf[25][11] ;
 wire \dp.rf.rf[25][12] ;
 wire \dp.rf.rf[25][13] ;
 wire \dp.rf.rf[25][14] ;
 wire \dp.rf.rf[25][15] ;
 wire \dp.rf.rf[25][16] ;
 wire \dp.rf.rf[25][17] ;
 wire \dp.rf.rf[25][18] ;
 wire \dp.rf.rf[25][19] ;
 wire \dp.rf.rf[25][1] ;
 wire \dp.rf.rf[25][20] ;
 wire \dp.rf.rf[25][21] ;
 wire \dp.rf.rf[25][22] ;
 wire \dp.rf.rf[25][23] ;
 wire \dp.rf.rf[25][24] ;
 wire \dp.rf.rf[25][25] ;
 wire \dp.rf.rf[25][26] ;
 wire \dp.rf.rf[25][27] ;
 wire \dp.rf.rf[25][28] ;
 wire \dp.rf.rf[25][29] ;
 wire \dp.rf.rf[25][2] ;
 wire \dp.rf.rf[25][30] ;
 wire \dp.rf.rf[25][31] ;
 wire \dp.rf.rf[25][3] ;
 wire \dp.rf.rf[25][4] ;
 wire \dp.rf.rf[25][5] ;
 wire \dp.rf.rf[25][6] ;
 wire \dp.rf.rf[25][7] ;
 wire \dp.rf.rf[25][8] ;
 wire \dp.rf.rf[25][9] ;
 wire \dp.rf.rf[26][0] ;
 wire \dp.rf.rf[26][10] ;
 wire \dp.rf.rf[26][11] ;
 wire \dp.rf.rf[26][12] ;
 wire \dp.rf.rf[26][13] ;
 wire \dp.rf.rf[26][14] ;
 wire \dp.rf.rf[26][15] ;
 wire \dp.rf.rf[26][16] ;
 wire \dp.rf.rf[26][17] ;
 wire \dp.rf.rf[26][18] ;
 wire \dp.rf.rf[26][19] ;
 wire \dp.rf.rf[26][1] ;
 wire \dp.rf.rf[26][20] ;
 wire \dp.rf.rf[26][21] ;
 wire \dp.rf.rf[26][22] ;
 wire \dp.rf.rf[26][23] ;
 wire \dp.rf.rf[26][24] ;
 wire \dp.rf.rf[26][25] ;
 wire \dp.rf.rf[26][26] ;
 wire \dp.rf.rf[26][27] ;
 wire \dp.rf.rf[26][28] ;
 wire \dp.rf.rf[26][29] ;
 wire \dp.rf.rf[26][2] ;
 wire \dp.rf.rf[26][30] ;
 wire \dp.rf.rf[26][31] ;
 wire \dp.rf.rf[26][3] ;
 wire \dp.rf.rf[26][4] ;
 wire \dp.rf.rf[26][5] ;
 wire \dp.rf.rf[26][6] ;
 wire \dp.rf.rf[26][7] ;
 wire \dp.rf.rf[26][8] ;
 wire \dp.rf.rf[26][9] ;
 wire \dp.rf.rf[27][0] ;
 wire \dp.rf.rf[27][10] ;
 wire \dp.rf.rf[27][11] ;
 wire \dp.rf.rf[27][12] ;
 wire \dp.rf.rf[27][13] ;
 wire \dp.rf.rf[27][14] ;
 wire \dp.rf.rf[27][15] ;
 wire \dp.rf.rf[27][16] ;
 wire \dp.rf.rf[27][17] ;
 wire \dp.rf.rf[27][18] ;
 wire \dp.rf.rf[27][19] ;
 wire \dp.rf.rf[27][1] ;
 wire \dp.rf.rf[27][20] ;
 wire \dp.rf.rf[27][21] ;
 wire \dp.rf.rf[27][22] ;
 wire \dp.rf.rf[27][23] ;
 wire \dp.rf.rf[27][24] ;
 wire \dp.rf.rf[27][25] ;
 wire \dp.rf.rf[27][26] ;
 wire \dp.rf.rf[27][27] ;
 wire \dp.rf.rf[27][28] ;
 wire \dp.rf.rf[27][29] ;
 wire \dp.rf.rf[27][2] ;
 wire \dp.rf.rf[27][30] ;
 wire \dp.rf.rf[27][31] ;
 wire \dp.rf.rf[27][3] ;
 wire \dp.rf.rf[27][4] ;
 wire \dp.rf.rf[27][5] ;
 wire \dp.rf.rf[27][6] ;
 wire \dp.rf.rf[27][7] ;
 wire \dp.rf.rf[27][8] ;
 wire \dp.rf.rf[27][9] ;
 wire \dp.rf.rf[28][0] ;
 wire \dp.rf.rf[28][10] ;
 wire \dp.rf.rf[28][11] ;
 wire \dp.rf.rf[28][12] ;
 wire \dp.rf.rf[28][13] ;
 wire \dp.rf.rf[28][14] ;
 wire \dp.rf.rf[28][15] ;
 wire \dp.rf.rf[28][16] ;
 wire \dp.rf.rf[28][17] ;
 wire \dp.rf.rf[28][18] ;
 wire \dp.rf.rf[28][19] ;
 wire \dp.rf.rf[28][1] ;
 wire \dp.rf.rf[28][20] ;
 wire \dp.rf.rf[28][21] ;
 wire \dp.rf.rf[28][22] ;
 wire \dp.rf.rf[28][23] ;
 wire \dp.rf.rf[28][24] ;
 wire \dp.rf.rf[28][25] ;
 wire \dp.rf.rf[28][26] ;
 wire \dp.rf.rf[28][27] ;
 wire \dp.rf.rf[28][28] ;
 wire \dp.rf.rf[28][29] ;
 wire \dp.rf.rf[28][2] ;
 wire \dp.rf.rf[28][30] ;
 wire \dp.rf.rf[28][31] ;
 wire \dp.rf.rf[28][3] ;
 wire \dp.rf.rf[28][4] ;
 wire \dp.rf.rf[28][5] ;
 wire \dp.rf.rf[28][6] ;
 wire \dp.rf.rf[28][7] ;
 wire \dp.rf.rf[28][8] ;
 wire \dp.rf.rf[28][9] ;
 wire \dp.rf.rf[29][0] ;
 wire \dp.rf.rf[29][10] ;
 wire \dp.rf.rf[29][11] ;
 wire \dp.rf.rf[29][12] ;
 wire \dp.rf.rf[29][13] ;
 wire \dp.rf.rf[29][14] ;
 wire \dp.rf.rf[29][15] ;
 wire \dp.rf.rf[29][16] ;
 wire \dp.rf.rf[29][17] ;
 wire \dp.rf.rf[29][18] ;
 wire \dp.rf.rf[29][19] ;
 wire \dp.rf.rf[29][1] ;
 wire \dp.rf.rf[29][20] ;
 wire \dp.rf.rf[29][21] ;
 wire \dp.rf.rf[29][22] ;
 wire \dp.rf.rf[29][23] ;
 wire \dp.rf.rf[29][24] ;
 wire \dp.rf.rf[29][25] ;
 wire \dp.rf.rf[29][26] ;
 wire \dp.rf.rf[29][27] ;
 wire \dp.rf.rf[29][28] ;
 wire \dp.rf.rf[29][29] ;
 wire \dp.rf.rf[29][2] ;
 wire \dp.rf.rf[29][30] ;
 wire \dp.rf.rf[29][31] ;
 wire \dp.rf.rf[29][3] ;
 wire \dp.rf.rf[29][4] ;
 wire \dp.rf.rf[29][5] ;
 wire \dp.rf.rf[29][6] ;
 wire \dp.rf.rf[29][7] ;
 wire \dp.rf.rf[29][8] ;
 wire \dp.rf.rf[29][9] ;
 wire \dp.rf.rf[2][0] ;
 wire \dp.rf.rf[2][10] ;
 wire \dp.rf.rf[2][11] ;
 wire \dp.rf.rf[2][12] ;
 wire \dp.rf.rf[2][13] ;
 wire \dp.rf.rf[2][14] ;
 wire \dp.rf.rf[2][15] ;
 wire \dp.rf.rf[2][16] ;
 wire \dp.rf.rf[2][17] ;
 wire \dp.rf.rf[2][18] ;
 wire \dp.rf.rf[2][19] ;
 wire \dp.rf.rf[2][1] ;
 wire \dp.rf.rf[2][20] ;
 wire \dp.rf.rf[2][21] ;
 wire \dp.rf.rf[2][22] ;
 wire \dp.rf.rf[2][23] ;
 wire \dp.rf.rf[2][24] ;
 wire \dp.rf.rf[2][25] ;
 wire \dp.rf.rf[2][26] ;
 wire \dp.rf.rf[2][27] ;
 wire \dp.rf.rf[2][28] ;
 wire \dp.rf.rf[2][29] ;
 wire \dp.rf.rf[2][2] ;
 wire \dp.rf.rf[2][30] ;
 wire \dp.rf.rf[2][31] ;
 wire \dp.rf.rf[2][3] ;
 wire \dp.rf.rf[2][4] ;
 wire \dp.rf.rf[2][5] ;
 wire \dp.rf.rf[2][6] ;
 wire \dp.rf.rf[2][7] ;
 wire \dp.rf.rf[2][8] ;
 wire \dp.rf.rf[2][9] ;
 wire \dp.rf.rf[30][0] ;
 wire \dp.rf.rf[30][10] ;
 wire \dp.rf.rf[30][11] ;
 wire \dp.rf.rf[30][12] ;
 wire \dp.rf.rf[30][13] ;
 wire \dp.rf.rf[30][14] ;
 wire \dp.rf.rf[30][15] ;
 wire \dp.rf.rf[30][16] ;
 wire \dp.rf.rf[30][17] ;
 wire \dp.rf.rf[30][18] ;
 wire \dp.rf.rf[30][19] ;
 wire \dp.rf.rf[30][1] ;
 wire \dp.rf.rf[30][20] ;
 wire \dp.rf.rf[30][21] ;
 wire \dp.rf.rf[30][22] ;
 wire \dp.rf.rf[30][23] ;
 wire \dp.rf.rf[30][24] ;
 wire \dp.rf.rf[30][25] ;
 wire \dp.rf.rf[30][26] ;
 wire \dp.rf.rf[30][27] ;
 wire \dp.rf.rf[30][28] ;
 wire \dp.rf.rf[30][29] ;
 wire \dp.rf.rf[30][2] ;
 wire \dp.rf.rf[30][30] ;
 wire \dp.rf.rf[30][31] ;
 wire \dp.rf.rf[30][3] ;
 wire \dp.rf.rf[30][4] ;
 wire \dp.rf.rf[30][5] ;
 wire \dp.rf.rf[30][6] ;
 wire \dp.rf.rf[30][7] ;
 wire \dp.rf.rf[30][8] ;
 wire \dp.rf.rf[30][9] ;
 wire \dp.rf.rf[31][0] ;
 wire \dp.rf.rf[31][10] ;
 wire \dp.rf.rf[31][11] ;
 wire \dp.rf.rf[31][12] ;
 wire \dp.rf.rf[31][13] ;
 wire \dp.rf.rf[31][14] ;
 wire \dp.rf.rf[31][15] ;
 wire \dp.rf.rf[31][16] ;
 wire \dp.rf.rf[31][17] ;
 wire \dp.rf.rf[31][18] ;
 wire \dp.rf.rf[31][19] ;
 wire \dp.rf.rf[31][1] ;
 wire \dp.rf.rf[31][20] ;
 wire \dp.rf.rf[31][21] ;
 wire \dp.rf.rf[31][22] ;
 wire \dp.rf.rf[31][23] ;
 wire \dp.rf.rf[31][24] ;
 wire \dp.rf.rf[31][25] ;
 wire \dp.rf.rf[31][26] ;
 wire \dp.rf.rf[31][27] ;
 wire \dp.rf.rf[31][28] ;
 wire \dp.rf.rf[31][29] ;
 wire \dp.rf.rf[31][2] ;
 wire \dp.rf.rf[31][30] ;
 wire \dp.rf.rf[31][31] ;
 wire \dp.rf.rf[31][3] ;
 wire \dp.rf.rf[31][4] ;
 wire \dp.rf.rf[31][5] ;
 wire \dp.rf.rf[31][6] ;
 wire \dp.rf.rf[31][7] ;
 wire \dp.rf.rf[31][8] ;
 wire \dp.rf.rf[31][9] ;
 wire \dp.rf.rf[3][0] ;
 wire \dp.rf.rf[3][10] ;
 wire \dp.rf.rf[3][11] ;
 wire \dp.rf.rf[3][12] ;
 wire \dp.rf.rf[3][13] ;
 wire \dp.rf.rf[3][14] ;
 wire \dp.rf.rf[3][15] ;
 wire \dp.rf.rf[3][16] ;
 wire \dp.rf.rf[3][17] ;
 wire \dp.rf.rf[3][18] ;
 wire \dp.rf.rf[3][19] ;
 wire \dp.rf.rf[3][1] ;
 wire \dp.rf.rf[3][20] ;
 wire \dp.rf.rf[3][21] ;
 wire \dp.rf.rf[3][22] ;
 wire \dp.rf.rf[3][23] ;
 wire \dp.rf.rf[3][24] ;
 wire \dp.rf.rf[3][25] ;
 wire \dp.rf.rf[3][26] ;
 wire \dp.rf.rf[3][27] ;
 wire \dp.rf.rf[3][28] ;
 wire \dp.rf.rf[3][29] ;
 wire \dp.rf.rf[3][2] ;
 wire \dp.rf.rf[3][30] ;
 wire \dp.rf.rf[3][31] ;
 wire \dp.rf.rf[3][3] ;
 wire \dp.rf.rf[3][4] ;
 wire \dp.rf.rf[3][5] ;
 wire \dp.rf.rf[3][6] ;
 wire \dp.rf.rf[3][7] ;
 wire \dp.rf.rf[3][8] ;
 wire \dp.rf.rf[3][9] ;
 wire \dp.rf.rf[4][0] ;
 wire \dp.rf.rf[4][10] ;
 wire \dp.rf.rf[4][11] ;
 wire \dp.rf.rf[4][12] ;
 wire \dp.rf.rf[4][13] ;
 wire \dp.rf.rf[4][14] ;
 wire \dp.rf.rf[4][15] ;
 wire \dp.rf.rf[4][16] ;
 wire \dp.rf.rf[4][17] ;
 wire \dp.rf.rf[4][18] ;
 wire \dp.rf.rf[4][19] ;
 wire \dp.rf.rf[4][1] ;
 wire \dp.rf.rf[4][20] ;
 wire \dp.rf.rf[4][21] ;
 wire \dp.rf.rf[4][22] ;
 wire \dp.rf.rf[4][23] ;
 wire \dp.rf.rf[4][24] ;
 wire \dp.rf.rf[4][25] ;
 wire \dp.rf.rf[4][26] ;
 wire \dp.rf.rf[4][27] ;
 wire \dp.rf.rf[4][28] ;
 wire \dp.rf.rf[4][29] ;
 wire \dp.rf.rf[4][2] ;
 wire \dp.rf.rf[4][30] ;
 wire \dp.rf.rf[4][31] ;
 wire \dp.rf.rf[4][3] ;
 wire \dp.rf.rf[4][4] ;
 wire \dp.rf.rf[4][5] ;
 wire \dp.rf.rf[4][6] ;
 wire \dp.rf.rf[4][7] ;
 wire \dp.rf.rf[4][8] ;
 wire \dp.rf.rf[4][9] ;
 wire \dp.rf.rf[5][0] ;
 wire \dp.rf.rf[5][10] ;
 wire \dp.rf.rf[5][11] ;
 wire \dp.rf.rf[5][12] ;
 wire \dp.rf.rf[5][13] ;
 wire \dp.rf.rf[5][14] ;
 wire \dp.rf.rf[5][15] ;
 wire \dp.rf.rf[5][16] ;
 wire \dp.rf.rf[5][17] ;
 wire \dp.rf.rf[5][18] ;
 wire \dp.rf.rf[5][19] ;
 wire \dp.rf.rf[5][1] ;
 wire \dp.rf.rf[5][20] ;
 wire \dp.rf.rf[5][21] ;
 wire \dp.rf.rf[5][22] ;
 wire \dp.rf.rf[5][23] ;
 wire \dp.rf.rf[5][24] ;
 wire \dp.rf.rf[5][25] ;
 wire \dp.rf.rf[5][26] ;
 wire \dp.rf.rf[5][27] ;
 wire \dp.rf.rf[5][28] ;
 wire \dp.rf.rf[5][29] ;
 wire \dp.rf.rf[5][2] ;
 wire \dp.rf.rf[5][30] ;
 wire \dp.rf.rf[5][31] ;
 wire \dp.rf.rf[5][3] ;
 wire \dp.rf.rf[5][4] ;
 wire \dp.rf.rf[5][5] ;
 wire \dp.rf.rf[5][6] ;
 wire \dp.rf.rf[5][7] ;
 wire \dp.rf.rf[5][8] ;
 wire \dp.rf.rf[5][9] ;
 wire \dp.rf.rf[6][0] ;
 wire \dp.rf.rf[6][10] ;
 wire \dp.rf.rf[6][11] ;
 wire \dp.rf.rf[6][12] ;
 wire \dp.rf.rf[6][13] ;
 wire \dp.rf.rf[6][14] ;
 wire \dp.rf.rf[6][15] ;
 wire \dp.rf.rf[6][16] ;
 wire \dp.rf.rf[6][17] ;
 wire \dp.rf.rf[6][18] ;
 wire \dp.rf.rf[6][19] ;
 wire \dp.rf.rf[6][1] ;
 wire \dp.rf.rf[6][20] ;
 wire \dp.rf.rf[6][21] ;
 wire \dp.rf.rf[6][22] ;
 wire \dp.rf.rf[6][23] ;
 wire \dp.rf.rf[6][24] ;
 wire \dp.rf.rf[6][25] ;
 wire \dp.rf.rf[6][26] ;
 wire \dp.rf.rf[6][27] ;
 wire \dp.rf.rf[6][28] ;
 wire \dp.rf.rf[6][29] ;
 wire \dp.rf.rf[6][2] ;
 wire \dp.rf.rf[6][30] ;
 wire \dp.rf.rf[6][31] ;
 wire \dp.rf.rf[6][3] ;
 wire \dp.rf.rf[6][4] ;
 wire \dp.rf.rf[6][5] ;
 wire \dp.rf.rf[6][6] ;
 wire \dp.rf.rf[6][7] ;
 wire \dp.rf.rf[6][8] ;
 wire \dp.rf.rf[6][9] ;
 wire \dp.rf.rf[7][0] ;
 wire \dp.rf.rf[7][10] ;
 wire \dp.rf.rf[7][11] ;
 wire \dp.rf.rf[7][12] ;
 wire \dp.rf.rf[7][13] ;
 wire \dp.rf.rf[7][14] ;
 wire \dp.rf.rf[7][15] ;
 wire \dp.rf.rf[7][16] ;
 wire \dp.rf.rf[7][17] ;
 wire \dp.rf.rf[7][18] ;
 wire \dp.rf.rf[7][19] ;
 wire \dp.rf.rf[7][1] ;
 wire \dp.rf.rf[7][20] ;
 wire \dp.rf.rf[7][21] ;
 wire \dp.rf.rf[7][22] ;
 wire \dp.rf.rf[7][23] ;
 wire \dp.rf.rf[7][24] ;
 wire \dp.rf.rf[7][25] ;
 wire \dp.rf.rf[7][26] ;
 wire \dp.rf.rf[7][27] ;
 wire \dp.rf.rf[7][28] ;
 wire \dp.rf.rf[7][29] ;
 wire \dp.rf.rf[7][2] ;
 wire \dp.rf.rf[7][30] ;
 wire \dp.rf.rf[7][31] ;
 wire \dp.rf.rf[7][3] ;
 wire \dp.rf.rf[7][4] ;
 wire \dp.rf.rf[7][5] ;
 wire \dp.rf.rf[7][6] ;
 wire \dp.rf.rf[7][7] ;
 wire \dp.rf.rf[7][8] ;
 wire \dp.rf.rf[7][9] ;
 wire \dp.rf.rf[8][0] ;
 wire \dp.rf.rf[8][10] ;
 wire \dp.rf.rf[8][11] ;
 wire \dp.rf.rf[8][12] ;
 wire \dp.rf.rf[8][13] ;
 wire \dp.rf.rf[8][14] ;
 wire \dp.rf.rf[8][15] ;
 wire \dp.rf.rf[8][16] ;
 wire \dp.rf.rf[8][17] ;
 wire \dp.rf.rf[8][18] ;
 wire \dp.rf.rf[8][19] ;
 wire \dp.rf.rf[8][1] ;
 wire \dp.rf.rf[8][20] ;
 wire \dp.rf.rf[8][21] ;
 wire \dp.rf.rf[8][22] ;
 wire \dp.rf.rf[8][23] ;
 wire \dp.rf.rf[8][24] ;
 wire \dp.rf.rf[8][25] ;
 wire \dp.rf.rf[8][26] ;
 wire \dp.rf.rf[8][27] ;
 wire \dp.rf.rf[8][28] ;
 wire \dp.rf.rf[8][29] ;
 wire \dp.rf.rf[8][2] ;
 wire \dp.rf.rf[8][30] ;
 wire \dp.rf.rf[8][31] ;
 wire \dp.rf.rf[8][3] ;
 wire \dp.rf.rf[8][4] ;
 wire \dp.rf.rf[8][5] ;
 wire \dp.rf.rf[8][6] ;
 wire \dp.rf.rf[8][7] ;
 wire \dp.rf.rf[8][8] ;
 wire \dp.rf.rf[8][9] ;
 wire \dp.rf.rf[9][0] ;
 wire \dp.rf.rf[9][10] ;
 wire \dp.rf.rf[9][11] ;
 wire \dp.rf.rf[9][12] ;
 wire \dp.rf.rf[9][13] ;
 wire \dp.rf.rf[9][14] ;
 wire \dp.rf.rf[9][15] ;
 wire \dp.rf.rf[9][16] ;
 wire \dp.rf.rf[9][17] ;
 wire \dp.rf.rf[9][18] ;
 wire \dp.rf.rf[9][19] ;
 wire \dp.rf.rf[9][1] ;
 wire \dp.rf.rf[9][20] ;
 wire \dp.rf.rf[9][21] ;
 wire \dp.rf.rf[9][22] ;
 wire \dp.rf.rf[9][23] ;
 wire \dp.rf.rf[9][24] ;
 wire \dp.rf.rf[9][25] ;
 wire \dp.rf.rf[9][26] ;
 wire \dp.rf.rf[9][27] ;
 wire \dp.rf.rf[9][28] ;
 wire \dp.rf.rf[9][29] ;
 wire \dp.rf.rf[9][2] ;
 wire \dp.rf.rf[9][30] ;
 wire \dp.rf.rf[9][31] ;
 wire \dp.rf.rf[9][3] ;
 wire \dp.rf.rf[9][4] ;
 wire \dp.rf.rf[9][5] ;
 wire \dp.rf.rf[9][6] ;
 wire \dp.rf.rf[9][7] ;
 wire \dp.rf.rf[9][8] ;
 wire \dp.rf.rf[9][9] ;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_buf_2 fanout1163 (.A(net1164),
    .X(net1163));
 sg13g2_inv_1 _08520_ (.Y(_02559_),
    .A(net1248));
 sg13g2_buf_2 fanout1162 (.A(net1204),
    .X(net1162));
 sg13g2_nor2b_2 _08522_ (.A(net27),
    .B_N(net1249),
    .Y(_02561_));
 sg13g2_buf_4 fanout1161 (.X(net1161),
    .A(net1162));
 sg13g2_buf_4 fanout1160 (.X(net1160),
    .A(net1161));
 sg13g2_buf_1 fanout1159 (.A(net1204),
    .X(net1159));
 sg13g2_and2_1 _08526_ (.A(net1),
    .B(net12),
    .X(_02565_));
 sg13g2_buf_4 fanout1158 (.X(net1158),
    .A(net1159));
 sg13g2_buf_4 fanout1157 (.X(net1157),
    .A(net1158));
 sg13g2_buf_2 fanout1156 (.A(net1157),
    .X(net1156));
 sg13g2_buf_4 fanout1155 (.X(net1155),
    .A(net1159));
 sg13g2_nor2_2 _08531_ (.A(net1251),
    .B(net1254),
    .Y(_02570_));
 sg13g2_buf_1 fanout1154 (.A(net1155),
    .X(net1154));
 sg13g2_nand4_1 _08533_ (.B(_02561_),
    .C(_02565_),
    .A(_02559_),
    .Y(_02572_),
    .D(_02570_));
 sg13g2_buf_2 fanout1153 (.A(net1155),
    .X(net1153));
 sg13g2_inv_4 _08535_ (.A(_02572_),
    .Y(net99));
 sg13g2_buf_1 fanout1152 (.A(net1159),
    .X(net1152));
 sg13g2_buf_4 fanout1151 (.X(net1151),
    .A(net1159));
 sg13g2_nor2_2 _08538_ (.A(net1243),
    .B(net1241),
    .Y(_02576_));
 sg13g2_buf_4 fanout1150 (.X(net1150),
    .A(net1152));
 sg13g2_and2_2 _08540_ (.A(net99),
    .B(_02576_),
    .X(_02578_));
 sg13g2_buf_2 fanout1149 (.A(net1204),
    .X(net1149));
 sg13g2_buf_1 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_1 fanout1147 (.A(net1148),
    .X(net1147));
 sg13g2_buf_4 fanout1146 (.X(net1146),
    .A(net1147));
 sg13g2_or2_1 _08545_ (.X(_02583_),
    .B(net1275),
    .A(net1258));
 sg13g2_buf_2 fanout1145 (.A(net1147),
    .X(net1145));
 sg13g2_buf_2 fanout1144 (.A(net1147),
    .X(net1144));
 sg13g2_buf_2 fanout1143 (.A(net1148),
    .X(net1143));
 sg13g2_buf_2 fanout1142 (.A(net1143),
    .X(net1142));
 sg13g2_buf_2 fanout1141 (.A(net1149),
    .X(net1141));
 sg13g2_buf_2 fanout1140 (.A(net1141),
    .X(net1140));
 sg13g2_buf_2 fanout1139 (.A(net1140),
    .X(net1139));
 sg13g2_buf_4 fanout1138 (.X(net1138),
    .A(net1141));
 sg13g2_nor3_2 _08554_ (.A(net1301),
    .B(net1342),
    .C(net1273),
    .Y(_02592_));
 sg13g2_nor2_1 _08555_ (.A(net1103),
    .B(_02592_),
    .Y(_02593_));
 sg13g2_buf_2 fanout1137 (.A(net1138),
    .X(net1137));
 sg13g2_buf_4 fanout1136 (.X(net1136),
    .A(net1141));
 sg13g2_buf_2 fanout1135 (.A(net1136),
    .X(net1135));
 sg13g2_mux4_1 _08559_ (.S0(net1357),
    .A0(\dp.rf.rf[2][8] ),
    .A1(\dp.rf.rf[3][8] ),
    .A2(\dp.rf.rf[10][8] ),
    .A3(\dp.rf.rf[11][8] ),
    .S1(net1273),
    .X(_02597_));
 sg13g2_mux4_1 _08560_ (.S0(net1357),
    .A0(\dp.rf.rf[0][8] ),
    .A1(\dp.rf.rf[1][8] ),
    .A2(\dp.rf.rf[8][8] ),
    .A3(\dp.rf.rf[9][8] ),
    .S1(net1269),
    .X(_02598_));
 sg13g2_buf_2 fanout1134 (.A(net1149),
    .X(net1134));
 sg13g2_buf_2 fanout1133 (.A(net1134),
    .X(net1133));
 sg13g2_inv_2 _08563_ (.Y(_02601_),
    .A(net1288));
 sg13g2_mux2_1 _08564_ (.A0(_02597_),
    .A1(_02598_),
    .S(net1101),
    .X(_02602_));
 sg13g2_nand2_1 _08565_ (.Y(_02603_),
    .A(_02593_),
    .B(_02602_));
 sg13g2_buf_4 fanout1132 (.X(net1132),
    .A(net1134));
 sg13g2_nand2_1 _08567_ (.Y(_02605_),
    .A(net1293),
    .B(net1266));
 sg13g2_buf_1 fanout1131 (.A(net1149),
    .X(net1131));
 sg13g2_buf_4 fanout1130 (.X(net1130),
    .A(net1131));
 sg13g2_buf_2 fanout1129 (.A(net1131),
    .X(net1129));
 sg13g2_nor2b_1 _08571_ (.A(net1374),
    .B_N(\dp.rf.rf[26][8] ),
    .Y(_02609_));
 sg13g2_a22oi_1 _08572_ (.Y(_02610_),
    .B1(net1098),
    .B2(_02609_),
    .A2(\dp.rf.rf[27][8] ),
    .A1(net1373));
 sg13g2_nand2b_1 _08573_ (.Y(_02611_),
    .B(net1266),
    .A_N(net1293));
 sg13g2_buf_2 fanout1128 (.A(net1129),
    .X(net1128));
 sg13g2_buf_4 fanout1127 (.X(net1127),
    .A(net1149));
 sg13g2_buf_4 fanout1126 (.X(net1126),
    .A(net1127));
 sg13g2_nor2b_1 _08577_ (.A(net1374),
    .B_N(\dp.rf.rf[24][8] ),
    .Y(_02615_));
 sg13g2_a22oi_1 _08578_ (.Y(_02616_),
    .B1(net1093),
    .B2(_02615_),
    .A2(\dp.rf.rf[25][8] ),
    .A1(net1373));
 sg13g2_buf_2 fanout1125 (.A(net1126),
    .X(net1125));
 sg13g2_buf_4 fanout1124 (.X(net1124),
    .A(net1127));
 sg13g2_buf_1 fanout1123 (.A(net9),
    .X(net1123));
 sg13g2_or2_1 _08582_ (.X(_02620_),
    .B(net1269),
    .A(net1292));
 sg13g2_buf_2 fanout1122 (.A(net1123),
    .X(net1122));
 sg13g2_buf_1 fanout1121 (.A(net1123),
    .X(net1121));
 sg13g2_buf_2 fanout1120 (.A(net1121),
    .X(net1120));
 sg13g2_nor2b_1 _08586_ (.A(net1373),
    .B_N(\dp.rf.rf[16][8] ),
    .Y(_02624_));
 sg13g2_a22oi_1 _08587_ (.Y(_02625_),
    .B1(net1084),
    .B2(_02624_),
    .A2(\dp.rf.rf[17][8] ),
    .A1(net1373));
 sg13g2_nand2b_1 _08588_ (.Y(_02626_),
    .B(net1294),
    .A_N(net1266));
 sg13g2_buf_1 fanout1119 (.A(net1121),
    .X(net1119));
 sg13g2_buf_1 fanout1118 (.A(net1119),
    .X(net1118));
 sg13g2_buf_2 fanout1117 (.A(net1119),
    .X(net1117));
 sg13g2_mux2_1 _08592_ (.A0(\dp.rf.rf[18][8] ),
    .A1(\dp.rf.rf[19][8] ),
    .S(net1373),
    .X(_02630_));
 sg13g2_nor2b_1 _08593_ (.A(net1275),
    .B_N(net1258),
    .Y(_02631_));
 sg13g2_buf_2 fanout1116 (.A(net1123),
    .X(net1116));
 sg13g2_o21ai_1 _08595_ (.B1(net1071),
    .Y(_02633_),
    .A1(net1077),
    .A2(_02630_));
 sg13g2_or4_1 _08596_ (.A(_02610_),
    .B(_02616_),
    .C(_02625_),
    .D(_02633_),
    .X(_02634_));
 sg13g2_nor2b_1 _08597_ (.A(net1282),
    .B_N(net1264),
    .Y(_02635_));
 sg13g2_buf_2 fanout1115 (.A(net1116),
    .X(net1115));
 sg13g2_nor2b_1 _08599_ (.A(net1258),
    .B_N(net1275),
    .Y(_02637_));
 sg13g2_buf_2 fanout1114 (.A(net1115),
    .X(net1114));
 sg13g2_buf_2 fanout1113 (.A(net1116),
    .X(net1113));
 sg13g2_mux2_1 _08602_ (.A0(\dp.rf.rf[12][8] ),
    .A1(\dp.rf.rf[13][8] ),
    .S(net1357),
    .X(_02640_));
 sg13g2_nand3_1 _08603_ (.B(net1064),
    .C(_02640_),
    .A(net1068),
    .Y(_02641_));
 sg13g2_and2_2 _08604_ (.A(net1284),
    .B(net1264),
    .X(_02642_));
 sg13g2_buf_2 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_buf_1 fanout1111 (.A(net1123),
    .X(net1111));
 sg13g2_mux2_1 _08607_ (.A0(\dp.rf.rf[14][8] ),
    .A1(\dp.rf.rf[15][8] ),
    .S(net1357),
    .X(_02645_));
 sg13g2_nand3_1 _08608_ (.B(net1063),
    .C(_02645_),
    .A(_02642_),
    .Y(_02646_));
 sg13g2_nor2_1 _08609_ (.A(net1282),
    .B(net1264),
    .Y(_02647_));
 sg13g2_buf_2 fanout1110 (.A(net1111),
    .X(net1110));
 sg13g2_and2_1 _08611_ (.A(net1260),
    .B(net1277),
    .X(_02649_));
 sg13g2_buf_2 fanout1109 (.A(net1111),
    .X(net1109));
 sg13g2_buf_2 fanout1108 (.A(net1109),
    .X(net1108));
 sg13g2_mux2_1 _08614_ (.A0(\dp.rf.rf[20][8] ),
    .A1(\dp.rf.rf[21][8] ),
    .S(net1357),
    .X(_02652_));
 sg13g2_nand3_1 _08615_ (.B(net1057),
    .C(_02652_),
    .A(net1060),
    .Y(_02653_));
 sg13g2_nor2b_1 _08616_ (.A(net1264),
    .B_N(net1284),
    .Y(_02654_));
 sg13g2_buf_2 fanout1107 (.A(net1109),
    .X(net1107));
 sg13g2_mux2_1 _08618_ (.A0(\dp.rf.rf[22][8] ),
    .A1(\dp.rf.rf[23][8] ),
    .S(net1373),
    .X(_02656_));
 sg13g2_nand3_1 _08619_ (.B(net1057),
    .C(_02656_),
    .A(net1053),
    .Y(_02657_));
 sg13g2_and4_1 _08620_ (.A(_02641_),
    .B(_02646_),
    .C(_02653_),
    .D(_02657_),
    .X(_02658_));
 sg13g2_mux2_1 _08621_ (.A0(\dp.rf.rf[4][8] ),
    .A1(\dp.rf.rf[5][8] ),
    .S(net1373),
    .X(_02659_));
 sg13g2_nand3_1 _08622_ (.B(net1064),
    .C(_02659_),
    .A(net1059),
    .Y(_02660_));
 sg13g2_mux2_1 _08623_ (.A0(\dp.rf.rf[6][8] ),
    .A1(\dp.rf.rf[7][8] ),
    .S(net1373),
    .X(_02661_));
 sg13g2_nand3_1 _08624_ (.B(net1064),
    .C(_02661_),
    .A(net1052),
    .Y(_02662_));
 sg13g2_and4_2 _08625_ (.A(net1258),
    .B(net1290),
    .C(net1275),
    .D(net1265),
    .X(_02663_));
 sg13g2_buf_2 fanout1106 (.A(net1109),
    .X(net1106));
 sg13g2_mux2_1 _08627_ (.A0(\dp.rf.rf[30][8] ),
    .A1(\dp.rf.rf[31][8] ),
    .S(net1374),
    .X(_02665_));
 sg13g2_nand2_1 _08628_ (.Y(_02666_),
    .A(_02663_),
    .B(_02665_));
 sg13g2_mux2_1 _08629_ (.A0(\dp.rf.rf[28][8] ),
    .A1(\dp.rf.rf[29][8] ),
    .S(net1374),
    .X(_02667_));
 sg13g2_nand3_1 _08630_ (.B(net1057),
    .C(_02667_),
    .A(net1068),
    .Y(_02668_));
 sg13g2_and4_1 _08631_ (.A(_02660_),
    .B(_02662_),
    .C(_02666_),
    .D(_02668_),
    .X(_02669_));
 sg13g2_and4_1 _08632_ (.A(_02603_),
    .B(_02634_),
    .C(_02658_),
    .D(_02669_),
    .X(_02670_));
 sg13g2_buf_2 fanout1105 (.A(_02583_),
    .X(net1105));
 sg13g2_nor2_1 _08634_ (.A(_02578_),
    .B(_02670_),
    .Y(net163));
 sg13g2_buf_1 fanout1104 (.A(net1105),
    .X(net1104));
 sg13g2_mux4_1 _08636_ (.S0(net1353),
    .A0(\dp.rf.rf[2][9] ),
    .A1(\dp.rf.rf[3][9] ),
    .A2(\dp.rf.rf[10][9] ),
    .A3(\dp.rf.rf[11][9] ),
    .S1(net1269),
    .X(_02673_));
 sg13g2_nor2_1 _08637_ (.A(net1101),
    .B(_02673_),
    .Y(_02674_));
 sg13g2_buf_2 fanout1103 (.A(net1105),
    .X(net1103));
 sg13g2_buf_2 fanout1102 (.A(_02601_),
    .X(net1102));
 sg13g2_a21oi_1 _08640_ (.A1(net1353),
    .A2(\dp.rf.rf[1][9] ),
    .Y(_02677_),
    .B1(net1082));
 sg13g2_buf_4 fanout1101 (.X(net1101),
    .A(_02601_));
 sg13g2_buf_2 fanout1100 (.A(_02605_),
    .X(net1100));
 sg13g2_buf_2 fanout1099 (.A(net1100),
    .X(net1099));
 sg13g2_buf_4 fanout1098 (.X(net1098),
    .A(net1099));
 sg13g2_buf_4 fanout1097 (.X(net1097),
    .A(net1099));
 sg13g2_nor2b_1 _08646_ (.A(net1353),
    .B_N(\dp.rf.rf[8][9] ),
    .Y(_02683_));
 sg13g2_a22oi_1 _08647_ (.Y(_02684_),
    .B1(net1090),
    .B2(_02683_),
    .A2(\dp.rf.rf[9][9] ),
    .A1(net1353));
 sg13g2_nor4_1 _08648_ (.A(net1103),
    .B(_02674_),
    .C(_02677_),
    .D(_02684_),
    .Y(_02685_));
 sg13g2_buf_4 fanout1096 (.X(net1096),
    .A(net1100));
 sg13g2_buf_4 fanout1095 (.X(net1095),
    .A(net1096));
 sg13g2_buf_1 fanout1094 (.A(_02611_),
    .X(net1094));
 sg13g2_buf_1 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_nor2b_1 _08653_ (.A(net1346),
    .B_N(\dp.rf.rf[26][9] ),
    .Y(_02690_));
 sg13g2_a22oi_1 _08654_ (.Y(_02691_),
    .B1(net1097),
    .B2(_02690_),
    .A2(\dp.rf.rf[27][9] ),
    .A1(net1346));
 sg13g2_nor2b_1 _08655_ (.A(net1346),
    .B_N(\dp.rf.rf[24][9] ),
    .Y(_02692_));
 sg13g2_a22oi_1 _08656_ (.Y(_02693_),
    .B1(net1090),
    .B2(_02692_),
    .A2(\dp.rf.rf[25][9] ),
    .A1(net1347));
 sg13g2_buf_2 fanout1092 (.A(net1093),
    .X(net1092));
 sg13g2_nor2b_1 _08658_ (.A(net1347),
    .B_N(\dp.rf.rf[16][9] ),
    .Y(_02695_));
 sg13g2_a22oi_1 _08659_ (.Y(_02696_),
    .B1(net1082),
    .B2(_02695_),
    .A2(\dp.rf.rf[17][9] ),
    .A1(net1347));
 sg13g2_buf_1 fanout1091 (.A(net1094),
    .X(net1091));
 sg13g2_buf_2 fanout1090 (.A(net1094),
    .X(net1090));
 sg13g2_mux2_1 _08662_ (.A0(\dp.rf.rf[18][9] ),
    .A1(\dp.rf.rf[19][9] ),
    .S(net1352),
    .X(_02699_));
 sg13g2_buf_1 fanout1089 (.A(net1094),
    .X(net1089));
 sg13g2_o21ai_1 _08664_ (.B1(net1070),
    .Y(_02701_),
    .A1(net1076),
    .A2(_02699_));
 sg13g2_nor4_1 _08665_ (.A(_02691_),
    .B(_02693_),
    .C(_02696_),
    .D(_02701_),
    .Y(_02702_));
 sg13g2_buf_2 fanout1088 (.A(net1089),
    .X(net1088));
 sg13g2_buf_1 fanout1087 (.A(net1089),
    .X(net1087));
 sg13g2_mux2_1 _08668_ (.A0(\dp.rf.rf[12][9] ),
    .A1(\dp.rf.rf[13][9] ),
    .S(net1349),
    .X(_02705_));
 sg13g2_nand3_1 _08669_ (.B(net1065),
    .C(_02705_),
    .A(net1067),
    .Y(_02706_));
 sg13g2_mux2_1 _08670_ (.A0(\dp.rf.rf[14][9] ),
    .A1(\dp.rf.rf[15][9] ),
    .S(net1349),
    .X(_02707_));
 sg13g2_nand3_1 _08671_ (.B(net1065),
    .C(_02707_),
    .A(_02642_),
    .Y(_02708_));
 sg13g2_buf_2 fanout1086 (.A(net1089),
    .X(net1086));
 sg13g2_buf_2 fanout1085 (.A(_02620_),
    .X(net1085));
 sg13g2_mux2_1 _08674_ (.A0(\dp.rf.rf[20][9] ),
    .A1(\dp.rf.rf[21][9] ),
    .S(net1347),
    .X(_02711_));
 sg13g2_nand3_1 _08675_ (.B(net1055),
    .C(_02711_),
    .A(net1059),
    .Y(_02712_));
 sg13g2_buf_4 fanout1084 (.X(net1084),
    .A(net1085));
 sg13g2_mux2_1 _08677_ (.A0(\dp.rf.rf[22][9] ),
    .A1(\dp.rf.rf[23][9] ),
    .S(net1347),
    .X(_02714_));
 sg13g2_nand3_1 _08678_ (.B(net1056),
    .C(_02714_),
    .A(net1052),
    .Y(_02715_));
 sg13g2_nand4_1 _08679_ (.B(_02708_),
    .C(_02712_),
    .A(_02706_),
    .Y(_02716_),
    .D(_02715_));
 sg13g2_buf_2 fanout1083 (.A(net1085),
    .X(net1083));
 sg13g2_mux2_1 _08681_ (.A0(\dp.rf.rf[4][9] ),
    .A1(\dp.rf.rf[5][9] ),
    .S(net1358),
    .X(_02718_));
 sg13g2_nand3_1 _08682_ (.B(net1065),
    .C(_02718_),
    .A(net1059),
    .Y(_02719_));
 sg13g2_mux2_1 _08683_ (.A0(\dp.rf.rf[6][9] ),
    .A1(\dp.rf.rf[7][9] ),
    .S(net1358),
    .X(_02720_));
 sg13g2_nand3_1 _08684_ (.B(net1065),
    .C(_02720_),
    .A(net1052),
    .Y(_02721_));
 sg13g2_buf_2 fanout1082 (.A(net1085),
    .X(net1082));
 sg13g2_buf_4 fanout1081 (.X(net1081),
    .A(_02620_));
 sg13g2_mux2_1 _08687_ (.A0(\dp.rf.rf[30][9] ),
    .A1(\dp.rf.rf[31][9] ),
    .S(net1349),
    .X(_02724_));
 sg13g2_nand2_1 _08688_ (.Y(_02725_),
    .A(_02663_),
    .B(_02724_));
 sg13g2_mux2_1 _08689_ (.A0(\dp.rf.rf[28][9] ),
    .A1(\dp.rf.rf[29][9] ),
    .S(net1353),
    .X(_02726_));
 sg13g2_nand3_1 _08690_ (.B(net1056),
    .C(_02726_),
    .A(_02635_),
    .Y(_02727_));
 sg13g2_nand4_1 _08691_ (.B(_02721_),
    .C(_02725_),
    .A(_02719_),
    .Y(_02728_),
    .D(_02727_));
 sg13g2_nor4_2 _08692_ (.A(_02685_),
    .B(_02702_),
    .C(_02716_),
    .Y(_02729_),
    .D(_02728_));
 sg13g2_nor2_1 _08693_ (.A(_02578_),
    .B(_02729_),
    .Y(net164));
 sg13g2_mux2_1 _08694_ (.A0(\dp.rf.rf[1][10] ),
    .A1(\dp.rf.rf[9][10] ),
    .S(net1268),
    .X(_02730_));
 sg13g2_nor2b_2 _08695_ (.A(net1332),
    .B_N(net1265),
    .Y(_02731_));
 sg13g2_buf_2 fanout1080 (.A(net1081),
    .X(net1080));
 sg13g2_buf_2 fanout1079 (.A(net1081),
    .X(net1079));
 sg13g2_buf_2 fanout1078 (.A(_02626_),
    .X(net1078));
 sg13g2_a221oi_1 _08699_ (.B2(\dp.rf.rf[8][10] ),
    .C1(net1295),
    .B1(_02731_),
    .A1(net1365),
    .Y(_02735_),
    .A2(_02730_));
 sg13g2_buf_2 fanout1077 (.A(net1078),
    .X(net1077));
 sg13g2_mux4_1 _08701_ (.S0(net1365),
    .A0(\dp.rf.rf[2][10] ),
    .A1(\dp.rf.rf[3][10] ),
    .A2(\dp.rf.rf[10][10] ),
    .A3(\dp.rf.rf[11][10] ),
    .S1(net1271),
    .X(_02737_));
 sg13g2_nor2_1 _08702_ (.A(net1258),
    .B(net1276),
    .Y(_02738_));
 sg13g2_buf_2 fanout1076 (.A(net1078),
    .X(net1076));
 sg13g2_buf_4 fanout1075 (.X(net1075),
    .A(_02626_));
 sg13g2_o21ai_1 _08705_ (.B1(net1051),
    .Y(_02741_),
    .A1(net1102),
    .A2(_02737_));
 sg13g2_or2_1 _08706_ (.X(_02742_),
    .B(_02741_),
    .A(_02735_));
 sg13g2_buf_2 fanout1074 (.A(net1075),
    .X(net1074));
 sg13g2_buf_4 fanout1073 (.X(net1073),
    .A(net1075));
 sg13g2_mux4_1 _08709_ (.S0(net1367),
    .A0(\dp.rf.rf[4][10] ),
    .A1(\dp.rf.rf[5][10] ),
    .A2(\dp.rf.rf[6][10] ),
    .A3(\dp.rf.rf[7][10] ),
    .S1(net1295),
    .X(_02745_));
 sg13g2_nand2b_2 _08710_ (.Y(_02746_),
    .B(net1276),
    .A_N(net1259));
 sg13g2_buf_2 fanout1072 (.A(_02631_),
    .X(net1072));
 sg13g2_nor2_2 _08712_ (.A(net1266),
    .B(_02746_),
    .Y(_02748_));
 sg13g2_buf_2 fanout1071 (.A(net1072),
    .X(net1071));
 sg13g2_buf_2 fanout1070 (.A(net1072),
    .X(net1070));
 sg13g2_buf_2 fanout1069 (.A(net1072),
    .X(net1069));
 sg13g2_mux4_1 _08716_ (.S0(net1365),
    .A0(\dp.rf.rf[12][10] ),
    .A1(\dp.rf.rf[13][10] ),
    .A2(\dp.rf.rf[14][10] ),
    .A3(\dp.rf.rf[15][10] ),
    .S1(net1295),
    .X(_02752_));
 sg13g2_and3_1 _08717_ (.X(_02753_),
    .A(net1268),
    .B(net1064),
    .C(_02752_));
 sg13g2_a21oi_1 _08718_ (.A1(_02745_),
    .A2(_02748_),
    .Y(_02754_),
    .B1(_02753_));
 sg13g2_buf_2 fanout1068 (.A(_02635_),
    .X(net1068));
 sg13g2_buf_2 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_1 fanout1066 (.A(_02637_),
    .X(net1066));
 sg13g2_nor2b_1 _08722_ (.A(net1378),
    .B_N(\dp.rf.rf[26][10] ),
    .Y(_02758_));
 sg13g2_a22oi_1 _08723_ (.Y(_02759_),
    .B1(net1099),
    .B2(_02758_),
    .A2(\dp.rf.rf[27][10] ),
    .A1(net1378));
 sg13g2_buf_2 fanout1065 (.A(net1066),
    .X(net1065));
 sg13g2_nor2b_1 _08725_ (.A(net1366),
    .B_N(\dp.rf.rf[16][10] ),
    .Y(_02761_));
 sg13g2_a22oi_1 _08726_ (.Y(_02762_),
    .B1(net1084),
    .B2(_02761_),
    .A2(\dp.rf.rf[17][10] ),
    .A1(net1366));
 sg13g2_nor2b_1 _08727_ (.A(net1378),
    .B_N(\dp.rf.rf[24][10] ),
    .Y(_02763_));
 sg13g2_a22oi_1 _08728_ (.Y(_02764_),
    .B1(net1092),
    .B2(_02763_),
    .A2(\dp.rf.rf[25][10] ),
    .A1(net1378));
 sg13g2_mux2_1 _08729_ (.A0(\dp.rf.rf[18][10] ),
    .A1(\dp.rf.rf[19][10] ),
    .S(net1366),
    .X(_02765_));
 sg13g2_o21ai_1 _08730_ (.B1(net1070),
    .Y(_02766_),
    .A1(net1077),
    .A2(_02765_));
 sg13g2_or4_1 _08731_ (.A(_02759_),
    .B(_02762_),
    .C(_02764_),
    .D(_02766_),
    .X(_02767_));
 sg13g2_nand2_2 _08732_ (.Y(_02768_),
    .A(net1258),
    .B(net1275));
 sg13g2_buf_2 fanout1064 (.A(net1065),
    .X(net1064));
 sg13g2_nor2_1 _08734_ (.A(net1267),
    .B(_02768_),
    .Y(_02770_));
 sg13g2_buf_2 fanout1063 (.A(net1066),
    .X(net1063));
 sg13g2_buf_1 fanout1062 (.A(net1066),
    .X(net1062));
 sg13g2_buf_2 fanout1061 (.A(net1066),
    .X(net1061));
 sg13g2_mux4_1 _08738_ (.S0(net1379),
    .A0(\dp.rf.rf[20][10] ),
    .A1(\dp.rf.rf[21][10] ),
    .A2(\dp.rf.rf[22][10] ),
    .A3(\dp.rf.rf[23][10] ),
    .S1(net1297),
    .X(_02774_));
 sg13g2_buf_2 fanout1060 (.A(_02647_),
    .X(net1060));
 sg13g2_mux2_1 _08740_ (.A0(\dp.rf.rf[30][10] ),
    .A1(\dp.rf.rf[31][10] ),
    .S(net1379),
    .X(_02776_));
 sg13g2_nand2_1 _08741_ (.Y(_02777_),
    .A(net1378),
    .B(\dp.rf.rf[29][10] ));
 sg13g2_nand2b_1 _08742_ (.Y(_02778_),
    .B(\dp.rf.rf[28][10] ),
    .A_N(net1378));
 sg13g2_a22oi_1 _08743_ (.Y(_02779_),
    .B1(net1092),
    .B2(_02768_),
    .A2(_02778_),
    .A1(_02777_));
 sg13g2_a221oi_1 _08744_ (.B2(_02663_),
    .C1(_02779_),
    .B1(_02776_),
    .A1(net952),
    .Y(_02780_),
    .A2(_02774_));
 sg13g2_nand4_1 _08745_ (.B(_02754_),
    .C(_02767_),
    .A(_02742_),
    .Y(_02781_),
    .D(_02780_));
 sg13g2_buf_2 fanout1059 (.A(net1060),
    .X(net1059));
 sg13g2_nor2b_1 _08747_ (.A(_02578_),
    .B_N(_02781_),
    .Y(net134));
 sg13g2_buf_1 fanout1058 (.A(_02649_),
    .X(net1058));
 sg13g2_buf_2 fanout1057 (.A(net1058),
    .X(net1057));
 sg13g2_nor2b_1 _08750_ (.A(net1382),
    .B_N(\dp.rf.rf[26][11] ),
    .Y(_02785_));
 sg13g2_a22oi_1 _08751_ (.Y(_02786_),
    .B1(net1098),
    .B2(_02785_),
    .A2(\dp.rf.rf[27][11] ),
    .A1(net1382));
 sg13g2_buf_2 fanout1056 (.A(net1057),
    .X(net1056));
 sg13g2_nor2b_1 _08753_ (.A(net1384),
    .B_N(\dp.rf.rf[16][11] ),
    .Y(_02788_));
 sg13g2_a22oi_1 _08754_ (.Y(_02789_),
    .B1(net1085),
    .B2(_02788_),
    .A2(\dp.rf.rf[17][11] ),
    .A1(net1384));
 sg13g2_buf_2 fanout1055 (.A(net1058),
    .X(net1055));
 sg13g2_buf_2 fanout1054 (.A(net1055),
    .X(net1054));
 sg13g2_nor2b_1 _08757_ (.A(net1382),
    .B_N(\dp.rf.rf[24][11] ),
    .Y(_02792_));
 sg13g2_a22oi_1 _08758_ (.Y(_02793_),
    .B1(net1093),
    .B2(_02792_),
    .A2(\dp.rf.rf[25][11] ),
    .A1(net1382));
 sg13g2_buf_2 fanout1053 (.A(_02654_),
    .X(net1053));
 sg13g2_mux2_1 _08760_ (.A0(\dp.rf.rf[18][11] ),
    .A1(\dp.rf.rf[19][11] ),
    .S(net1385),
    .X(_02795_));
 sg13g2_buf_2 fanout1052 (.A(net1053),
    .X(net1052));
 sg13g2_o21ai_1 _08762_ (.B1(net1071),
    .Y(_02797_),
    .A1(net1077),
    .A2(_02795_));
 sg13g2_nor4_1 _08763_ (.A(_02786_),
    .B(_02789_),
    .C(_02793_),
    .D(_02797_),
    .Y(_02798_));
 sg13g2_mux2_1 _08764_ (.A0(\dp.rf.rf[1][11] ),
    .A1(\dp.rf.rf[9][11] ),
    .S(net1270),
    .X(_02799_));
 sg13g2_a221oi_1 _08765_ (.B2(net1377),
    .C1(net1297),
    .B1(_02799_),
    .A1(\dp.rf.rf[8][11] ),
    .Y(_02800_),
    .A2(_02731_));
 sg13g2_nand2b_1 _08766_ (.Y(_02801_),
    .B(net1297),
    .A_N(net1376));
 sg13g2_buf_2 fanout1051 (.A(_02738_),
    .X(net1051));
 sg13g2_nor2b_1 _08768_ (.A(net1270),
    .B_N(\dp.rf.rf[2][11] ),
    .Y(_02803_));
 sg13g2_a22oi_1 _08769_ (.Y(_02804_),
    .B1(_02801_),
    .B2(_02803_),
    .A2(\dp.rf.rf[10][11] ),
    .A1(net1270));
 sg13g2_nand2_1 _08770_ (.Y(_02805_),
    .A(net1297),
    .B(net1376));
 sg13g2_nor2b_1 _08771_ (.A(net1270),
    .B_N(\dp.rf.rf[3][11] ),
    .Y(_02806_));
 sg13g2_a22oi_1 _08772_ (.Y(_02807_),
    .B1(_02805_),
    .B2(_02806_),
    .A2(\dp.rf.rf[11][11] ),
    .A1(net1270));
 sg13g2_nor4_1 _08773_ (.A(net1103),
    .B(_02800_),
    .C(_02804_),
    .D(_02807_),
    .Y(_02808_));
 sg13g2_buf_4 fanout1050 (.X(net1050),
    .A(_02738_));
 sg13g2_mux4_1 _08775_ (.S0(net1386),
    .A0(\dp.rf.rf[20][11] ),
    .A1(\dp.rf.rf[21][11] ),
    .A2(\dp.rf.rf[22][11] ),
    .A3(\dp.rf.rf[23][11] ),
    .S1(net1299),
    .X(_02810_));
 sg13g2_mux4_1 _08776_ (.S0(net1380),
    .A0(\dp.rf.rf[28][11] ),
    .A1(\dp.rf.rf[29][11] ),
    .A2(\dp.rf.rf[30][11] ),
    .A3(\dp.rf.rf[31][11] ),
    .S1(net1297),
    .X(_02811_));
 sg13g2_and3_1 _08777_ (.X(_02812_),
    .A(net1272),
    .B(net1057),
    .C(_02811_));
 sg13g2_a21o_1 _08778_ (.A2(_02810_),
    .A1(net952),
    .B1(_02812_),
    .X(_02813_));
 sg13g2_mux4_1 _08779_ (.S0(net1388),
    .A0(\dp.rf.rf[4][11] ),
    .A1(\dp.rf.rf[5][11] ),
    .A2(\dp.rf.rf[6][11] ),
    .A3(\dp.rf.rf[7][11] ),
    .S1(net1299),
    .X(_02814_));
 sg13g2_nand3b_1 _08780_ (.B(net1277),
    .C(net1270),
    .Y(_02815_),
    .A_N(net1260));
 sg13g2_buf_1 fanout1049 (.A(_02856_),
    .X(net1049));
 sg13g2_mux4_1 _08782_ (.S0(net1377),
    .A0(\dp.rf.rf[12][11] ),
    .A1(\dp.rf.rf[13][11] ),
    .A2(\dp.rf.rf[14][11] ),
    .A3(\dp.rf.rf[15][11] ),
    .S1(net1297),
    .X(_02817_));
 sg13g2_nor2b_1 _08783_ (.A(_02815_),
    .B_N(_02817_),
    .Y(_02818_));
 sg13g2_a21o_1 _08784_ (.A2(_02814_),
    .A1(_02748_),
    .B1(_02818_),
    .X(_02819_));
 sg13g2_nor4_2 _08785_ (.A(_02798_),
    .B(_02808_),
    .C(_02813_),
    .Y(_02820_),
    .D(_02819_));
 sg13g2_nor2_1 _08786_ (.A(_02578_),
    .B(_02820_),
    .Y(net135));
 sg13g2_buf_4 fanout1048 (.X(net1048),
    .A(_02856_));
 sg13g2_nand4_1 _08788_ (.B(net1301),
    .C(net1277),
    .A(net1260),
    .Y(_02822_),
    .D(net1273));
 sg13g2_buf_2 fanout1047 (.A(_02856_),
    .X(net1047));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(net1047));
 sg13g2_buf_1 fanout1045 (.A(net1047),
    .X(net1045));
 sg13g2_nor2b_1 _08792_ (.A(net1368),
    .B_N(\dp.rf.rf[30][12] ),
    .Y(_02826_));
 sg13g2_a21oi_1 _08793_ (.A1(net1368),
    .A2(\dp.rf.rf[31][12] ),
    .Y(_02827_),
    .B1(_02826_));
 sg13g2_mux2_1 _08794_ (.A0(\dp.rf.rf[28][12] ),
    .A1(\dp.rf.rf[29][12] ),
    .S(net1368),
    .X(_02828_));
 sg13g2_nand3_1 _08795_ (.B(net1056),
    .C(_02828_),
    .A(net1068),
    .Y(_02829_));
 sg13g2_o21ai_1 _08796_ (.B1(_02829_),
    .Y(_02830_),
    .A1(_02822_),
    .A2(_02827_));
 sg13g2_nand2_1 _08797_ (.Y(_02831_),
    .A(net1367),
    .B(\dp.rf.rf[23][12] ));
 sg13g2_nand2b_1 _08798_ (.Y(_02832_),
    .B(\dp.rf.rf[22][12] ),
    .A_N(net1367));
 sg13g2_a22oi_1 _08799_ (.Y(_02833_),
    .B1(net1078),
    .B2(_02768_),
    .A2(_02832_),
    .A1(_02831_));
 sg13g2_nand2_1 _08800_ (.Y(_02834_),
    .A(net1367),
    .B(\dp.rf.rf[21][12] ));
 sg13g2_nand2b_1 _08801_ (.Y(_02835_),
    .B(\dp.rf.rf[20][12] ),
    .A_N(net1367));
 sg13g2_a22oi_1 _08802_ (.Y(_02836_),
    .B1(net1083),
    .B2(_02768_),
    .A2(_02835_),
    .A1(_02834_));
 sg13g2_buf_2 fanout1044 (.A(net1047),
    .X(net1044));
 sg13g2_buf_1 fanout1043 (.A(_02929_),
    .X(net1043));
 sg13g2_nor2b_1 _08805_ (.A(net1367),
    .B_N(\dp.rf.rf[26][12] ),
    .Y(_02839_));
 sg13g2_a22oi_1 _08806_ (.Y(_02840_),
    .B1(net1099),
    .B2(_02839_),
    .A2(\dp.rf.rf[27][12] ),
    .A1(net1366));
 sg13g2_nor2b_1 _08807_ (.A(net1366),
    .B_N(\dp.rf.rf[16][12] ),
    .Y(_02841_));
 sg13g2_a22oi_1 _08808_ (.Y(_02842_),
    .B1(net1083),
    .B2(_02841_),
    .A2(\dp.rf.rf[17][12] ),
    .A1(net1366));
 sg13g2_nor2b_1 _08809_ (.A(net1367),
    .B_N(\dp.rf.rf[24][12] ),
    .Y(_02843_));
 sg13g2_a22oi_1 _08810_ (.Y(_02844_),
    .B1(net1091),
    .B2(_02843_),
    .A2(\dp.rf.rf[25][12] ),
    .A1(net1366));
 sg13g2_mux2_1 _08811_ (.A0(\dp.rf.rf[18][12] ),
    .A1(\dp.rf.rf[19][12] ),
    .S(net1366),
    .X(_02845_));
 sg13g2_o21ai_1 _08812_ (.B1(net1070),
    .Y(_02846_),
    .A1(net1076),
    .A2(_02845_));
 sg13g2_nor4_1 _08813_ (.A(_02840_),
    .B(_02842_),
    .C(_02844_),
    .D(_02846_),
    .Y(_02847_));
 sg13g2_nor4_2 _08814_ (.A(_02830_),
    .B(_02833_),
    .C(_02836_),
    .Y(_02848_),
    .D(_02847_));
 sg13g2_buf_2 fanout1042 (.A(_02929_),
    .X(net1042));
 sg13g2_nand2_1 _08816_ (.Y(_02850_),
    .A(net1376),
    .B(\dp.rf.rf[1][12] ));
 sg13g2_buf_2 fanout1041 (.A(_03654_),
    .X(net1041));
 sg13g2_nor2b_1 _08818_ (.A(net1376),
    .B_N(\dp.rf.rf[8][12] ),
    .Y(_02852_));
 sg13g2_a22oi_1 _08819_ (.Y(_02853_),
    .B1(net1092),
    .B2(_02852_),
    .A2(\dp.rf.rf[9][12] ),
    .A1(net1376));
 sg13g2_buf_2 fanout1040 (.A(_03654_),
    .X(net1040));
 sg13g2_a22oi_1 _08821_ (.Y(_02855_),
    .B1(_02853_),
    .B2(net1104),
    .A2(_02850_),
    .A1(net1059));
 sg13g2_inv_2 _08822_ (.Y(_02856_),
    .A(net1262));
 sg13g2_buf_1 fanout1039 (.A(_03662_),
    .X(net1039));
 sg13g2_and2_1 _08824_ (.A(net1271),
    .B(\dp.rf.rf[11][12] ),
    .X(_02858_));
 sg13g2_a22oi_1 _08825_ (.Y(_02859_),
    .B1(_02805_),
    .B2(_02858_),
    .A2(\dp.rf.rf[3][12] ),
    .A1(net1049));
 sg13g2_buf_2 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_nor2b_1 _08827_ (.A(net1270),
    .B_N(\dp.rf.rf[2][12] ),
    .Y(_02861_));
 sg13g2_a22oi_1 _08828_ (.Y(_02862_),
    .B1(_02801_),
    .B2(_02861_),
    .A2(\dp.rf.rf[10][12] ),
    .A1(net1270));
 sg13g2_nor2_1 _08829_ (.A(_02859_),
    .B(_02862_),
    .Y(_02863_));
 sg13g2_nor2b_1 _08830_ (.A(net1376),
    .B_N(\dp.rf.rf[14][12] ),
    .Y(_02864_));
 sg13g2_a22oi_1 _08831_ (.Y(_02865_),
    .B1(net1099),
    .B2(_02864_),
    .A2(\dp.rf.rf[15][12] ),
    .A1(net1376));
 sg13g2_buf_2 fanout1037 (.A(net1038),
    .X(net1037));
 sg13g2_nor2b_1 _08833_ (.A(net1376),
    .B_N(\dp.rf.rf[12][12] ),
    .Y(_02867_));
 sg13g2_a22oi_1 _08834_ (.Y(_02868_),
    .B1(net1092),
    .B2(_02867_),
    .A2(\dp.rf.rf[13][12] ),
    .A1(net1377));
 sg13g2_buf_2 fanout1036 (.A(net1038),
    .X(net1036));
 sg13g2_nor2b_1 _08836_ (.A(net1379),
    .B_N(\dp.rf.rf[4][12] ),
    .Y(_02870_));
 sg13g2_a22oi_1 _08837_ (.Y(_02871_),
    .B1(net1084),
    .B2(_02870_),
    .A2(\dp.rf.rf[5][12] ),
    .A1(net1379));
 sg13g2_mux2_1 _08838_ (.A0(\dp.rf.rf[6][12] ),
    .A1(\dp.rf.rf[7][12] ),
    .S(net1379),
    .X(_02872_));
 sg13g2_o21ai_1 _08839_ (.B1(net1064),
    .Y(_02873_),
    .A1(net1077),
    .A2(_02872_));
 sg13g2_nor4_1 _08840_ (.A(_02865_),
    .B(_02868_),
    .C(_02871_),
    .D(_02873_),
    .Y(_02874_));
 sg13g2_a21oi_1 _08841_ (.A1(_02855_),
    .A2(_02863_),
    .Y(_02875_),
    .B1(_02874_));
 sg13g2_and2_1 _08842_ (.A(_02848_),
    .B(_02875_),
    .X(_02876_));
 sg13g2_buf_2 fanout1035 (.A(net1038),
    .X(net1035));
 sg13g2_nor2_1 _08844_ (.A(_02578_),
    .B(_02876_),
    .Y(net136));
 sg13g2_nor2b_1 _08845_ (.A(net1342),
    .B_N(\dp.rf.rf[30][13] ),
    .Y(_02878_));
 sg13g2_a21oi_1 _08846_ (.A1(net1342),
    .A2(\dp.rf.rf[31][13] ),
    .Y(_02879_),
    .B1(_02878_));
 sg13g2_mux2_1 _08847_ (.A0(\dp.rf.rf[28][13] ),
    .A1(\dp.rf.rf[29][13] ),
    .S(net1342),
    .X(_02880_));
 sg13g2_nand3_1 _08848_ (.B(net1058),
    .C(_02880_),
    .A(net1068),
    .Y(_02881_));
 sg13g2_o21ai_1 _08849_ (.B1(_02881_),
    .Y(_02882_),
    .A1(_02822_),
    .A2(_02879_));
 sg13g2_buf_2 fanout1034 (.A(net1035),
    .X(net1034));
 sg13g2_mux2_1 _08851_ (.A0(\dp.rf.rf[20][13] ),
    .A1(\dp.rf.rf[21][13] ),
    .S(net1371),
    .X(_02884_));
 sg13g2_nand3_1 _08852_ (.B(net1054),
    .C(_02884_),
    .A(net1060),
    .Y(_02885_));
 sg13g2_mux2_1 _08853_ (.A0(\dp.rf.rf[22][13] ),
    .A1(\dp.rf.rf[23][13] ),
    .S(net1371),
    .X(_02886_));
 sg13g2_nand3_1 _08854_ (.B(net1058),
    .C(_02886_),
    .A(net1052),
    .Y(_02887_));
 sg13g2_nand2_1 _08855_ (.Y(_02888_),
    .A(_02885_),
    .B(_02887_));
 sg13g2_mux2_1 _08856_ (.A0(\dp.rf.rf[12][13] ),
    .A1(\dp.rf.rf[13][13] ),
    .S(net1355),
    .X(_02889_));
 sg13g2_nand3_1 _08857_ (.B(net1063),
    .C(_02889_),
    .A(net1068),
    .Y(_02890_));
 sg13g2_mux2_1 _08858_ (.A0(\dp.rf.rf[14][13] ),
    .A1(\dp.rf.rf[15][13] ),
    .S(net1355),
    .X(_02891_));
 sg13g2_nand3_1 _08859_ (.B(net1063),
    .C(_02891_),
    .A(_02642_),
    .Y(_02892_));
 sg13g2_mux2_1 _08860_ (.A0(\dp.rf.rf[4][13] ),
    .A1(\dp.rf.rf[5][13] ),
    .S(net1372),
    .X(_02893_));
 sg13g2_nand3_1 _08861_ (.B(net1063),
    .C(_02893_),
    .A(_02647_),
    .Y(_02894_));
 sg13g2_mux2_1 _08862_ (.A0(\dp.rf.rf[6][13] ),
    .A1(\dp.rf.rf[7][13] ),
    .S(net1372),
    .X(_02895_));
 sg13g2_nand3_1 _08863_ (.B(net1063),
    .C(_02895_),
    .A(net1053),
    .Y(_02896_));
 sg13g2_nand4_1 _08864_ (.B(_02892_),
    .C(_02894_),
    .A(_02890_),
    .Y(_02897_),
    .D(_02896_));
 sg13g2_nor3_1 _08865_ (.A(_02882_),
    .B(_02888_),
    .C(_02897_),
    .Y(_02898_));
 sg13g2_buf_1 fanout1033 (.A(net1039),
    .X(net1033));
 sg13g2_mux4_1 _08867_ (.S0(net1359),
    .A0(\dp.rf.rf[8][13] ),
    .A1(\dp.rf.rf[9][13] ),
    .A2(\dp.rf.rf[10][13] ),
    .A3(\dp.rf.rf[11][13] ),
    .S1(net1291),
    .X(_02900_));
 sg13g2_buf_2 fanout1032 (.A(net1033),
    .X(net1032));
 sg13g2_nor2_1 _08869_ (.A(net1049),
    .B(net1104),
    .Y(_02902_));
 sg13g2_nor2b_1 _08870_ (.A(net1371),
    .B_N(\dp.rf.rf[18][13] ),
    .Y(_02903_));
 sg13g2_a22oi_1 _08871_ (.Y(_02904_),
    .B1(net1077),
    .B2(_02903_),
    .A2(\dp.rf.rf[19][13] ),
    .A1(net1371));
 sg13g2_nor2b_1 _08872_ (.A(net1371),
    .B_N(\dp.rf.rf[16][13] ),
    .Y(_02905_));
 sg13g2_a22oi_1 _08873_ (.Y(_02906_),
    .B1(net1084),
    .B2(_02905_),
    .A2(\dp.rf.rf[17][13] ),
    .A1(net1371));
 sg13g2_nor2b_1 _08874_ (.A(net1371),
    .B_N(\dp.rf.rf[26][13] ),
    .Y(_02907_));
 sg13g2_a22oi_1 _08875_ (.Y(_02908_),
    .B1(net1098),
    .B2(_02907_),
    .A2(\dp.rf.rf[27][13] ),
    .A1(net1371));
 sg13g2_nor2b_1 _08876_ (.A(net1342),
    .B_N(\dp.rf.rf[24][13] ),
    .Y(_02909_));
 sg13g2_a22oi_1 _08877_ (.Y(_02910_),
    .B1(net1089),
    .B2(_02909_),
    .A2(\dp.rf.rf[25][13] ),
    .A1(net1342));
 sg13g2_nor4_1 _08878_ (.A(_02904_),
    .B(_02906_),
    .C(_02908_),
    .D(_02910_),
    .Y(_02911_));
 sg13g2_mux2_1 _08879_ (.A0(\dp.rf.rf[2][13] ),
    .A1(\dp.rf.rf[3][13] ),
    .S(net1372),
    .X(_02912_));
 sg13g2_nand2_1 _08880_ (.Y(_02913_),
    .A(net1301),
    .B(_02912_));
 sg13g2_nand3_1 _08881_ (.B(net1372),
    .C(\dp.rf.rf[1][13] ),
    .A(net1102),
    .Y(_02914_));
 sg13g2_a22oi_1 _08882_ (.Y(_02915_),
    .B1(net1273),
    .B2(net1104),
    .A2(_02914_),
    .A1(_02913_));
 sg13g2_a221oi_1 _08883_ (.B2(net1071),
    .C1(_02915_),
    .B1(_02911_),
    .A1(_02900_),
    .Y(_02916_),
    .A2(_02902_));
 sg13g2_and2_1 _08884_ (.A(_02898_),
    .B(_02916_),
    .X(_02917_));
 sg13g2_buf_1 fanout1031 (.A(net1033),
    .X(net1031));
 sg13g2_nor2_1 _08886_ (.A(_02578_),
    .B(_02917_),
    .Y(net137));
 sg13g2_nor2b_1 _08887_ (.A(net1324),
    .B_N(\dp.rf.rf[18][14] ),
    .Y(_02919_));
 sg13g2_a22oi_1 _08888_ (.Y(_02920_),
    .B1(net1073),
    .B2(_02919_),
    .A2(\dp.rf.rf[19][14] ),
    .A1(net1324));
 sg13g2_nor2b_1 _08889_ (.A(net1324),
    .B_N(\dp.rf.rf[16][14] ),
    .Y(_02921_));
 sg13g2_a22oi_1 _08890_ (.Y(_02922_),
    .B1(net1079),
    .B2(_02921_),
    .A2(\dp.rf.rf[17][14] ),
    .A1(net1324));
 sg13g2_nor2b_1 _08891_ (.A(net1324),
    .B_N(\dp.rf.rf[26][14] ),
    .Y(_02923_));
 sg13g2_a22oi_1 _08892_ (.Y(_02924_),
    .B1(net1095),
    .B2(_02923_),
    .A2(\dp.rf.rf[27][14] ),
    .A1(net1324));
 sg13g2_mux2_1 _08893_ (.A0(\dp.rf.rf[24][14] ),
    .A1(\dp.rf.rf[25][14] ),
    .S(net1329),
    .X(_02925_));
 sg13g2_o21ai_1 _08894_ (.B1(net1069),
    .Y(_02926_),
    .A1(net1086),
    .A2(_02925_));
 sg13g2_or4_1 _08895_ (.A(_02920_),
    .B(_02922_),
    .C(_02924_),
    .D(_02926_),
    .X(_02927_));
 sg13g2_mux4_1 _08896_ (.S0(net1325),
    .A0(\dp.rf.rf[20][14] ),
    .A1(\dp.rf.rf[21][14] ),
    .A2(\dp.rf.rf[22][14] ),
    .A3(\dp.rf.rf[23][14] ),
    .S1(net1284),
    .X(_02928_));
 sg13g2_nand3_1 _08897_ (.B(net1275),
    .C(net1265),
    .A(net1258),
    .Y(_02929_));
 sg13g2_buf_2 fanout1030 (.A(net1033),
    .X(net1030));
 sg13g2_buf_1 fanout1029 (.A(net1039),
    .X(net1029));
 sg13g2_mux4_1 _08900_ (.S0(net1327),
    .A0(\dp.rf.rf[28][14] ),
    .A1(\dp.rf.rf[29][14] ),
    .A2(\dp.rf.rf[30][14] ),
    .A3(\dp.rf.rf[31][14] ),
    .S1(net1285),
    .X(_02932_));
 sg13g2_nor2b_1 _08901_ (.A(net1042),
    .B_N(_02932_),
    .Y(_02933_));
 sg13g2_a21oi_1 _08902_ (.A1(net951),
    .A2(_02928_),
    .Y(_02934_),
    .B1(_02933_));
 sg13g2_buf_2 fanout1028 (.A(net1029),
    .X(net1028));
 sg13g2_mux2_1 _08904_ (.A0(\dp.rf.rf[8][14] ),
    .A1(\dp.rf.rf[9][14] ),
    .S(net1325),
    .X(_02936_));
 sg13g2_mux2_1 _08905_ (.A0(\dp.rf.rf[10][14] ),
    .A1(\dp.rf.rf[11][14] ),
    .S(net1326),
    .X(_02937_));
 sg13g2_and2_1 _08906_ (.A(net1326),
    .B(\dp.rf.rf[1][14] ),
    .X(_02938_));
 sg13g2_mux2_1 _08907_ (.A0(\dp.rf.rf[2][14] ),
    .A1(\dp.rf.rf[3][14] ),
    .S(net1326),
    .X(_02939_));
 sg13g2_mux4_1 _08908_ (.S0(net1285),
    .A0(_02936_),
    .A1(_02937_),
    .A2(_02938_),
    .A3(_02939_),
    .S1(net1045),
    .X(_02940_));
 sg13g2_nand2_1 _08909_ (.Y(_02941_),
    .A(net1050),
    .B(_02940_));
 sg13g2_mux4_1 _08910_ (.S0(net1324),
    .A0(\dp.rf.rf[12][14] ),
    .A1(\dp.rf.rf[13][14] ),
    .A2(\dp.rf.rf[14][14] ),
    .A3(\dp.rf.rf[15][14] ),
    .S1(net1284),
    .X(_02942_));
 sg13g2_mux4_1 _08911_ (.S0(net1325),
    .A0(\dp.rf.rf[4][14] ),
    .A1(\dp.rf.rf[5][14] ),
    .A2(\dp.rf.rf[6][14] ),
    .A3(\dp.rf.rf[7][14] ),
    .S1(net1284),
    .X(_02943_));
 sg13g2_mux2_1 _08912_ (.A0(_02942_),
    .A1(_02943_),
    .S(net1045),
    .X(_02944_));
 sg13g2_nand2_1 _08913_ (.Y(_02945_),
    .A(net1062),
    .B(_02944_));
 sg13g2_and4_2 _08914_ (.A(_02927_),
    .B(_02934_),
    .C(_02941_),
    .D(_02945_),
    .X(_02946_));
 sg13g2_buf_1 fanout1027 (.A(net1029),
    .X(net1027));
 sg13g2_nor2_1 _08916_ (.A(_02578_),
    .B(_02946_),
    .Y(net138));
 sg13g2_mux4_1 _08917_ (.S0(net1351),
    .A0(\dp.rf.rf[20][15] ),
    .A1(\dp.rf.rf[21][15] ),
    .A2(\dp.rf.rf[22][15] ),
    .A3(\dp.rf.rf[23][15] ),
    .S1(net1293),
    .X(_02948_));
 sg13g2_mux4_1 _08918_ (.S0(net1360),
    .A0(\dp.rf.rf[28][15] ),
    .A1(\dp.rf.rf[29][15] ),
    .A2(\dp.rf.rf[30][15] ),
    .A3(\dp.rf.rf[31][15] ),
    .S1(net1293),
    .X(_02949_));
 sg13g2_nor2b_1 _08919_ (.A(net1043),
    .B_N(_02949_),
    .Y(_02950_));
 sg13g2_a21oi_1 _08920_ (.A1(net952),
    .A2(_02948_),
    .Y(_02951_),
    .B1(_02950_));
 sg13g2_mux4_1 _08921_ (.S0(net1361),
    .A0(\dp.rf.rf[2][15] ),
    .A1(\dp.rf.rf[3][15] ),
    .A2(\dp.rf.rf[10][15] ),
    .A3(\dp.rf.rf[11][15] ),
    .S1(net1266),
    .X(_02952_));
 sg13g2_mux4_1 _08922_ (.S0(net1353),
    .A0(\dp.rf.rf[0][15] ),
    .A1(\dp.rf.rf[1][15] ),
    .A2(\dp.rf.rf[8][15] ),
    .A3(\dp.rf.rf[9][15] ),
    .S1(net1266),
    .X(_02953_));
 sg13g2_mux2_1 _08923_ (.A0(_02952_),
    .A1(_02953_),
    .S(net1102),
    .X(_02954_));
 sg13g2_nand2_1 _08924_ (.Y(_02955_),
    .A(_02593_),
    .B(_02954_));
 sg13g2_nor2b_1 _08925_ (.A(net1351),
    .B_N(\dp.rf.rf[18][15] ),
    .Y(_02956_));
 sg13g2_a22oi_1 _08926_ (.Y(_02957_),
    .B1(net1076),
    .B2(_02956_),
    .A2(\dp.rf.rf[19][15] ),
    .A1(net1351));
 sg13g2_nor2b_1 _08927_ (.A(net1351),
    .B_N(\dp.rf.rf[16][15] ),
    .Y(_02958_));
 sg13g2_a22oi_1 _08928_ (.Y(_02959_),
    .B1(net1082),
    .B2(_02958_),
    .A2(\dp.rf.rf[17][15] ),
    .A1(net1351));
 sg13g2_nor2b_1 _08929_ (.A(net1351),
    .B_N(\dp.rf.rf[26][15] ),
    .Y(_02960_));
 sg13g2_a22oi_1 _08930_ (.Y(_02961_),
    .B1(net1097),
    .B2(_02960_),
    .A2(\dp.rf.rf[27][15] ),
    .A1(net1351));
 sg13g2_mux2_1 _08931_ (.A0(\dp.rf.rf[24][15] ),
    .A1(\dp.rf.rf[25][15] ),
    .S(net1351),
    .X(_02962_));
 sg13g2_o21ai_1 _08932_ (.B1(net1070),
    .Y(_02963_),
    .A1(net1090),
    .A2(_02962_));
 sg13g2_or4_1 _08933_ (.A(_02957_),
    .B(_02959_),
    .C(_02961_),
    .D(_02963_),
    .X(_02964_));
 sg13g2_nor2b_1 _08934_ (.A(net1361),
    .B_N(\dp.rf.rf[6][15] ),
    .Y(_02965_));
 sg13g2_a22oi_1 _08935_ (.Y(_02966_),
    .B1(net1076),
    .B2(_02965_),
    .A2(\dp.rf.rf[7][15] ),
    .A1(net1361));
 sg13g2_nor2b_1 _08936_ (.A(net1360),
    .B_N(\dp.rf.rf[4][15] ),
    .Y(_02967_));
 sg13g2_a22oi_1 _08937_ (.Y(_02968_),
    .B1(net1083),
    .B2(_02967_),
    .A2(\dp.rf.rf[5][15] ),
    .A1(net1360));
 sg13g2_nor2b_1 _08938_ (.A(net1360),
    .B_N(\dp.rf.rf[14][15] ),
    .Y(_02969_));
 sg13g2_a22oi_1 _08939_ (.Y(_02970_),
    .B1(net1099),
    .B2(_02969_),
    .A2(\dp.rf.rf[15][15] ),
    .A1(net1360));
 sg13g2_mux2_1 _08940_ (.A0(\dp.rf.rf[12][15] ),
    .A1(\dp.rf.rf[13][15] ),
    .S(net1360),
    .X(_02971_));
 sg13g2_o21ai_1 _08941_ (.B1(net1065),
    .Y(_02972_),
    .A1(net1091),
    .A2(_02971_));
 sg13g2_or4_1 _08942_ (.A(_02966_),
    .B(_02968_),
    .C(_02970_),
    .D(_02972_),
    .X(_02973_));
 sg13g2_and4_1 _08943_ (.A(_02951_),
    .B(_02955_),
    .C(_02964_),
    .D(_02973_),
    .X(_02974_));
 sg13g2_nor2_1 _08944_ (.A(_02578_),
    .B(_02974_),
    .Y(net139));
 sg13g2_buf_2 fanout1026 (.A(net1029),
    .X(net1026));
 sg13g2_nor2_1 _08946_ (.A(net1239),
    .B(_02572_),
    .Y(_02976_));
 sg13g2_buf_2 fanout1025 (.A(net1026),
    .X(net1025));
 sg13g2_nor2b_1 _08948_ (.A(net1352),
    .B_N(\dp.rf.rf[26][16] ),
    .Y(_02978_));
 sg13g2_a22oi_1 _08949_ (.Y(_02979_),
    .B1(net1097),
    .B2(_02978_),
    .A2(\dp.rf.rf[27][16] ),
    .A1(net1352));
 sg13g2_nor2b_1 _08950_ (.A(net1352),
    .B_N(\dp.rf.rf[24][16] ),
    .Y(_02980_));
 sg13g2_a22oi_1 _08951_ (.Y(_02981_),
    .B1(net1090),
    .B2(_02980_),
    .A2(\dp.rf.rf[25][16] ),
    .A1(net1352));
 sg13g2_nor2b_1 _08952_ (.A(net1352),
    .B_N(\dp.rf.rf[16][16] ),
    .Y(_02982_));
 sg13g2_a22oi_1 _08953_ (.Y(_02983_),
    .B1(net1082),
    .B2(_02982_),
    .A2(\dp.rf.rf[17][16] ),
    .A1(net1352));
 sg13g2_mux2_1 _08954_ (.A0(\dp.rf.rf[18][16] ),
    .A1(\dp.rf.rf[19][16] ),
    .S(net1352),
    .X(_02984_));
 sg13g2_o21ai_1 _08955_ (.B1(net1070),
    .Y(_02985_),
    .A1(net1076),
    .A2(_02984_));
 sg13g2_nor4_1 _08956_ (.A(_02979_),
    .B(_02981_),
    .C(_02983_),
    .D(_02985_),
    .Y(_02986_));
 sg13g2_mux2_1 _08957_ (.A0(\dp.rf.rf[20][16] ),
    .A1(\dp.rf.rf[21][16] ),
    .S(net1354),
    .X(_02987_));
 sg13g2_nand3_1 _08958_ (.B(net1056),
    .C(_02987_),
    .A(net1059),
    .Y(_02988_));
 sg13g2_mux2_1 _08959_ (.A0(\dp.rf.rf[30][16] ),
    .A1(\dp.rf.rf[31][16] ),
    .S(net1353),
    .X(_02989_));
 sg13g2_nand2_1 _08960_ (.Y(_02990_),
    .A(_02663_),
    .B(_02989_));
 sg13g2_mux2_1 _08961_ (.A0(\dp.rf.rf[22][16] ),
    .A1(\dp.rf.rf[23][16] ),
    .S(net1353),
    .X(_02991_));
 sg13g2_nand3_1 _08962_ (.B(net1056),
    .C(_02991_),
    .A(net1052),
    .Y(_02992_));
 sg13g2_mux2_1 _08963_ (.A0(\dp.rf.rf[28][16] ),
    .A1(\dp.rf.rf[29][16] ),
    .S(net1354),
    .X(_02993_));
 sg13g2_nand3_1 _08964_ (.B(net1056),
    .C(_02993_),
    .A(net1068),
    .Y(_02994_));
 sg13g2_nand4_1 _08965_ (.B(_02990_),
    .C(_02992_),
    .A(_02988_),
    .Y(_02995_),
    .D(_02994_));
 sg13g2_mux4_1 _08966_ (.S0(net1361),
    .A0(\dp.rf.rf[4][16] ),
    .A1(\dp.rf.rf[5][16] ),
    .A2(\dp.rf.rf[6][16] ),
    .A3(\dp.rf.rf[7][16] ),
    .S1(net1293),
    .X(_02996_));
 sg13g2_mux4_1 _08967_ (.S0(net1364),
    .A0(\dp.rf.rf[12][16] ),
    .A1(\dp.rf.rf[13][16] ),
    .A2(\dp.rf.rf[14][16] ),
    .A3(\dp.rf.rf[15][16] ),
    .S1(net1295),
    .X(_02997_));
 sg13g2_nor2b_1 _08968_ (.A(_02815_),
    .B_N(_02997_),
    .Y(_02998_));
 sg13g2_a21o_1 _08969_ (.A2(_02996_),
    .A1(_02748_),
    .B1(_02998_),
    .X(_02999_));
 sg13g2_buf_1 fanout1024 (.A(_03666_),
    .X(net1024));
 sg13g2_mux4_1 _08971_ (.S0(net1354),
    .A0(\dp.rf.rf[2][16] ),
    .A1(\dp.rf.rf[3][16] ),
    .A2(\dp.rf.rf[10][16] ),
    .A3(\dp.rf.rf[11][16] ),
    .S1(net1266),
    .X(_03001_));
 sg13g2_inv_1 _08972_ (.Y(_03002_),
    .A(_03001_));
 sg13g2_mux2_1 _08973_ (.A0(\dp.rf.rf[1][16] ),
    .A1(\dp.rf.rf[9][16] ),
    .S(net1266),
    .X(_03003_));
 sg13g2_buf_2 fanout1023 (.A(net1024),
    .X(net1023));
 sg13g2_a221oi_1 _08975_ (.B2(net1354),
    .C1(net1292),
    .B1(_03003_),
    .A1(\dp.rf.rf[8][16] ),
    .Y(_03005_),
    .A2(_02731_));
 sg13g2_a22oi_1 _08976_ (.Y(_03006_),
    .B1(_03005_),
    .B2(net1103),
    .A2(_03002_),
    .A1(net1292));
 sg13g2_nor4_2 _08977_ (.A(_02986_),
    .B(_02995_),
    .C(_02999_),
    .Y(_03007_),
    .D(_03006_));
 sg13g2_nor2_1 _08978_ (.A(_02976_),
    .B(_03007_),
    .Y(net140));
 sg13g2_buf_2 fanout1022 (.A(net1023),
    .X(net1022));
 sg13g2_nor2b_1 _08980_ (.A(net1340),
    .B_N(\dp.rf.rf[30][17] ),
    .Y(_03009_));
 sg13g2_a21oi_1 _08981_ (.A1(net1340),
    .A2(\dp.rf.rf[31][17] ),
    .Y(_03010_),
    .B1(_03009_));
 sg13g2_mux2_1 _08982_ (.A0(\dp.rf.rf[28][17] ),
    .A1(\dp.rf.rf[29][17] ),
    .S(net1340),
    .X(_03011_));
 sg13g2_nand3_1 _08983_ (.B(net1054),
    .C(_03011_),
    .A(net1067),
    .Y(_03012_));
 sg13g2_o21ai_1 _08984_ (.B1(_03012_),
    .Y(_03013_),
    .A1(_02822_),
    .A2(_03010_));
 sg13g2_mux2_1 _08985_ (.A0(\dp.rf.rf[22][17] ),
    .A1(\dp.rf.rf[23][17] ),
    .S(net1343),
    .X(_03014_));
 sg13g2_nand3_1 _08986_ (.B(net1054),
    .C(_03014_),
    .A(net1053),
    .Y(_03015_));
 sg13g2_mux2_1 _08987_ (.A0(\dp.rf.rf[20][17] ),
    .A1(\dp.rf.rf[21][17] ),
    .S(net1343),
    .X(_03016_));
 sg13g2_nand3_1 _08988_ (.B(net1054),
    .C(_03016_),
    .A(net1060),
    .Y(_03017_));
 sg13g2_nand2_1 _08989_ (.Y(_03018_),
    .A(_03015_),
    .B(_03017_));
 sg13g2_buf_2 fanout1021 (.A(net1023),
    .X(net1021));
 sg13g2_mux2_1 _08991_ (.A0(\dp.rf.rf[12][17] ),
    .A1(\dp.rf.rf[13][17] ),
    .S(net1340),
    .X(_03020_));
 sg13g2_nand3_1 _08992_ (.B(net1062),
    .C(_03020_),
    .A(net1067),
    .Y(_03021_));
 sg13g2_mux2_1 _08993_ (.A0(\dp.rf.rf[14][17] ),
    .A1(\dp.rf.rf[15][17] ),
    .S(net1327),
    .X(_03022_));
 sg13g2_nand3_1 _08994_ (.B(net1062),
    .C(_03022_),
    .A(_02642_),
    .Y(_03023_));
 sg13g2_mux2_1 _08995_ (.A0(\dp.rf.rf[4][17] ),
    .A1(\dp.rf.rf[5][17] ),
    .S(net1340),
    .X(_03024_));
 sg13g2_nand3_1 _08996_ (.B(net1062),
    .C(_03024_),
    .A(net1060),
    .Y(_03025_));
 sg13g2_mux2_1 _08997_ (.A0(\dp.rf.rf[6][17] ),
    .A1(\dp.rf.rf[7][17] ),
    .S(net1341),
    .X(_03026_));
 sg13g2_nand3_1 _08998_ (.B(net1061),
    .C(_03026_),
    .A(net1053),
    .Y(_03027_));
 sg13g2_nand4_1 _08999_ (.B(_03023_),
    .C(_03025_),
    .A(_03021_),
    .Y(_03028_),
    .D(_03027_));
 sg13g2_nor3_1 _09000_ (.A(_03013_),
    .B(_03018_),
    .C(_03028_),
    .Y(_03029_));
 sg13g2_buf_2 fanout1020 (.A(net1021),
    .X(net1020));
 sg13g2_nor2b_1 _09002_ (.A(net1341),
    .B_N(\dp.rf.rf[26][17] ),
    .Y(_03031_));
 sg13g2_a22oi_1 _09003_ (.Y(_03032_),
    .B1(net1096),
    .B2(_03031_),
    .A2(\dp.rf.rf[27][17] ),
    .A1(net1341));
 sg13g2_nor2b_1 _09004_ (.A(net1341),
    .B_N(\dp.rf.rf[24][17] ),
    .Y(_03033_));
 sg13g2_a22oi_1 _09005_ (.Y(_03034_),
    .B1(net1088),
    .B2(_03033_),
    .A2(\dp.rf.rf[25][17] ),
    .A1(net1341));
 sg13g2_nor2b_1 _09006_ (.A(net1341),
    .B_N(\dp.rf.rf[18][17] ),
    .Y(_03035_));
 sg13g2_a22oi_1 _09007_ (.Y(_03036_),
    .B1(net1075),
    .B2(_03035_),
    .A2(\dp.rf.rf[19][17] ),
    .A1(net1341));
 sg13g2_buf_1 fanout1019 (.A(net1024),
    .X(net1019));
 sg13g2_nor2b_1 _09009_ (.A(net1344),
    .B_N(\dp.rf.rf[16][17] ),
    .Y(_03038_));
 sg13g2_a22oi_1 _09010_ (.Y(_03039_),
    .B1(net1081),
    .B2(_03038_),
    .A2(\dp.rf.rf[17][17] ),
    .A1(net1344));
 sg13g2_nor4_1 _09011_ (.A(_03032_),
    .B(_03034_),
    .C(_03036_),
    .D(_03039_),
    .Y(_03040_));
 sg13g2_buf_2 fanout1018 (.A(net1019),
    .X(net1018));
 sg13g2_mux4_1 _09013_ (.S0(net1340),
    .A0(\dp.rf.rf[2][17] ),
    .A1(\dp.rf.rf[3][17] ),
    .A2(\dp.rf.rf[10][17] ),
    .A3(\dp.rf.rf[11][17] ),
    .S1(net1265),
    .X(_03042_));
 sg13g2_inv_1 _09014_ (.Y(_03043_),
    .A(_03042_));
 sg13g2_mux2_1 _09015_ (.A0(\dp.rf.rf[1][17] ),
    .A1(\dp.rf.rf[9][17] ),
    .S(net1274),
    .X(_03044_));
 sg13g2_buf_1 fanout1017 (.A(net1019),
    .X(net1017));
 sg13g2_a221oi_1 _09017_ (.B2(net1340),
    .C1(net1290),
    .B1(_03044_),
    .A1(\dp.rf.rf[8][17] ),
    .Y(_03046_),
    .A2(_02731_));
 sg13g2_a22oi_1 _09018_ (.Y(_03047_),
    .B1(_03046_),
    .B2(net1105),
    .A2(_03043_),
    .A1(net1290));
 sg13g2_a21oi_2 _09019_ (.B1(_03047_),
    .Y(_03048_),
    .A2(_03040_),
    .A1(net1072));
 sg13g2_a21oi_1 _09020_ (.A1(_03029_),
    .A2(_03048_),
    .Y(net141),
    .B1(_02976_));
 sg13g2_nand2_2 _09021_ (.Y(_03049_),
    .A(net1051),
    .B(_02592_));
 sg13g2_o21ai_1 _09022_ (.B1(_03049_),
    .Y(_03050_),
    .A1(net1239),
    .A2(_02572_));
 sg13g2_buf_2 fanout1016 (.A(net1019),
    .X(net1016));
 sg13g2_mux4_1 _09024_ (.S0(net1320),
    .A0(\dp.rf.rf[20][18] ),
    .A1(\dp.rf.rf[21][18] ),
    .A2(\dp.rf.rf[22][18] ),
    .A3(\dp.rf.rf[23][18] ),
    .S1(net1283),
    .X(_03052_));
 sg13g2_mux4_1 _09025_ (.S0(net1346),
    .A0(\dp.rf.rf[28][18] ),
    .A1(\dp.rf.rf[29][18] ),
    .A2(\dp.rf.rf[30][18] ),
    .A3(\dp.rf.rf[31][18] ),
    .S1(net1292),
    .X(_03053_));
 sg13g2_nor2b_1 _09026_ (.A(net1042),
    .B_N(_03053_),
    .Y(_03054_));
 sg13g2_a21o_1 _09027_ (.A2(_03052_),
    .A1(net951),
    .B1(_03054_),
    .X(_03055_));
 sg13g2_mux4_1 _09028_ (.S0(net1320),
    .A0(\dp.rf.rf[4][18] ),
    .A1(\dp.rf.rf[5][18] ),
    .A2(\dp.rf.rf[6][18] ),
    .A3(\dp.rf.rf[7][18] ),
    .S1(net1292),
    .X(_03056_));
 sg13g2_mux4_1 _09029_ (.S0(net1346),
    .A0(\dp.rf.rf[12][18] ),
    .A1(\dp.rf.rf[13][18] ),
    .A2(\dp.rf.rf[14][18] ),
    .A3(\dp.rf.rf[15][18] ),
    .S1(net1292),
    .X(_03057_));
 sg13g2_nor2b_1 _09030_ (.A(_02815_),
    .B_N(_03057_),
    .Y(_03058_));
 sg13g2_a21o_1 _09031_ (.A2(_03056_),
    .A1(_02748_),
    .B1(_03058_),
    .X(_03059_));
 sg13g2_nor2b_1 _09032_ (.A(net1346),
    .B_N(\dp.rf.rf[18][18] ),
    .Y(_03060_));
 sg13g2_a22oi_1 _09033_ (.Y(_03061_),
    .B1(net1076),
    .B2(_03060_),
    .A2(\dp.rf.rf[19][18] ),
    .A1(net1346));
 sg13g2_nor2b_1 _09034_ (.A(net1348),
    .B_N(\dp.rf.rf[16][18] ),
    .Y(_03062_));
 sg13g2_a22oi_1 _09035_ (.Y(_03063_),
    .B1(net1082),
    .B2(_03062_),
    .A2(\dp.rf.rf[17][18] ),
    .A1(net1348));
 sg13g2_nor2b_1 _09036_ (.A(net1320),
    .B_N(\dp.rf.rf[26][18] ),
    .Y(_03064_));
 sg13g2_a22oi_1 _09037_ (.Y(_03065_),
    .B1(net1097),
    .B2(_03064_),
    .A2(\dp.rf.rf[27][18] ),
    .A1(net1320));
 sg13g2_mux2_1 _09038_ (.A0(\dp.rf.rf[24][18] ),
    .A1(\dp.rf.rf[25][18] ),
    .S(net1346),
    .X(_03066_));
 sg13g2_o21ai_1 _09039_ (.B1(net1069),
    .Y(_03067_),
    .A1(net1090),
    .A2(_03066_));
 sg13g2_nor4_1 _09040_ (.A(_03061_),
    .B(_03063_),
    .C(_03065_),
    .D(_03067_),
    .Y(_03068_));
 sg13g2_nor2b_1 _09041_ (.A(net1348),
    .B_N(\dp.rf.rf[10][18] ),
    .Y(_03069_));
 sg13g2_a22oi_1 _09042_ (.Y(_03070_),
    .B1(net1097),
    .B2(_03069_),
    .A2(\dp.rf.rf[11][18] ),
    .A1(net1348));
 sg13g2_nor2b_1 _09043_ (.A(net1321),
    .B_N(\dp.rf.rf[8][18] ),
    .Y(_03071_));
 sg13g2_a22oi_1 _09044_ (.Y(_03072_),
    .B1(net1087),
    .B2(_03071_),
    .A2(\dp.rf.rf[9][18] ),
    .A1(net1348));
 sg13g2_nor2b_1 _09045_ (.A(net1348),
    .B_N(\dp.rf.rf[0][18] ),
    .Y(_03073_));
 sg13g2_a22oi_1 _09046_ (.Y(_03074_),
    .B1(net1082),
    .B2(_03073_),
    .A2(\dp.rf.rf[1][18] ),
    .A1(net1348));
 sg13g2_mux2_1 _09047_ (.A0(\dp.rf.rf[2][18] ),
    .A1(\dp.rf.rf[3][18] ),
    .S(net1348),
    .X(_03075_));
 sg13g2_o21ai_1 _09048_ (.B1(net1050),
    .Y(_03076_),
    .A1(net1076),
    .A2(_03075_));
 sg13g2_nor4_1 _09049_ (.A(_03070_),
    .B(_03072_),
    .C(_03074_),
    .D(_03076_),
    .Y(_03077_));
 sg13g2_nor4_2 _09050_ (.A(_03055_),
    .B(_03059_),
    .C(_03068_),
    .Y(_03078_),
    .D(_03077_));
 sg13g2_nor2_1 _09051_ (.A(_03050_),
    .B(_03078_),
    .Y(net142));
 sg13g2_mux4_1 _09052_ (.S0(net1326),
    .A0(\dp.rf.rf[4][19] ),
    .A1(\dp.rf.rf[5][19] ),
    .A2(\dp.rf.rf[6][19] ),
    .A3(\dp.rf.rf[7][19] ),
    .S1(net1285),
    .X(_03079_));
 sg13g2_nand2_1 _09053_ (.Y(_03080_),
    .A(_02748_),
    .B(_03079_));
 sg13g2_mux4_1 _09054_ (.S0(net1320),
    .A0(\dp.rf.rf[12][19] ),
    .A1(\dp.rf.rf[13][19] ),
    .A2(\dp.rf.rf[14][19] ),
    .A3(\dp.rf.rf[15][19] ),
    .S1(net1283),
    .X(_03081_));
 sg13g2_nand2_1 _09055_ (.Y(_03082_),
    .A(net1061),
    .B(_03081_));
 sg13g2_mux4_1 _09056_ (.S0(net1321),
    .A0(\dp.rf.rf[8][19] ),
    .A1(\dp.rf.rf[9][19] ),
    .A2(\dp.rf.rf[10][19] ),
    .A3(\dp.rf.rf[11][19] ),
    .S1(net1283),
    .X(_03083_));
 sg13g2_nand2_1 _09057_ (.Y(_03084_),
    .A(net1050),
    .B(_03083_));
 sg13g2_a21oi_1 _09058_ (.A1(_03082_),
    .A2(_03084_),
    .Y(_03085_),
    .B1(net1045));
 sg13g2_nor2b_1 _09059_ (.A(net1321),
    .B_N(\dp.rf.rf[26][19] ),
    .Y(_03086_));
 sg13g2_a22oi_1 _09060_ (.Y(_03087_),
    .B1(net1096),
    .B2(_03086_),
    .A2(\dp.rf.rf[27][19] ),
    .A1(net1321));
 sg13g2_nor2b_1 _09061_ (.A(net1321),
    .B_N(\dp.rf.rf[24][19] ),
    .Y(_03088_));
 sg13g2_a22oi_1 _09062_ (.Y(_03089_),
    .B1(net1087),
    .B2(_03088_),
    .A2(\dp.rf.rf[25][19] ),
    .A1(net1322));
 sg13g2_nor2b_1 _09063_ (.A(net1322),
    .B_N(\dp.rf.rf[16][19] ),
    .Y(_03090_));
 sg13g2_a22oi_1 _09064_ (.Y(_03091_),
    .B1(net1080),
    .B2(_03090_),
    .A2(\dp.rf.rf[17][19] ),
    .A1(net1322));
 sg13g2_mux2_1 _09065_ (.A0(\dp.rf.rf[18][19] ),
    .A1(\dp.rf.rf[19][19] ),
    .S(net1322),
    .X(_03092_));
 sg13g2_o21ai_1 _09066_ (.B1(net1069),
    .Y(_03093_),
    .A1(net1074),
    .A2(_03092_));
 sg13g2_nor4_1 _09067_ (.A(_03087_),
    .B(_03089_),
    .C(_03091_),
    .D(_03093_),
    .Y(_03094_));
 sg13g2_mux2_1 _09068_ (.A0(\dp.rf.rf[2][19] ),
    .A1(\dp.rf.rf[3][19] ),
    .S(net1326),
    .X(_03095_));
 sg13g2_nand2_1 _09069_ (.Y(_03096_),
    .A(net1291),
    .B(_03095_));
 sg13g2_nor2b_2 _09070_ (.A(net1291),
    .B_N(net1357),
    .Y(_03097_));
 sg13g2_nand2_1 _09071_ (.Y(_03098_),
    .A(\dp.rf.rf[1][19] ),
    .B(_03097_));
 sg13g2_a22oi_1 _09072_ (.Y(_03099_),
    .B1(net1269),
    .B2(net1103),
    .A2(_03098_),
    .A1(_03096_));
 sg13g2_mux2_1 _09073_ (.A0(\dp.rf.rf[30][19] ),
    .A1(\dp.rf.rf[31][19] ),
    .S(net1326),
    .X(_03100_));
 sg13g2_nand2_1 _09074_ (.Y(_03101_),
    .A(_02663_),
    .B(_03100_));
 sg13g2_mux2_1 _09075_ (.A0(\dp.rf.rf[22][19] ),
    .A1(\dp.rf.rf[23][19] ),
    .S(net1326),
    .X(_03102_));
 sg13g2_nand3_1 _09076_ (.B(net1055),
    .C(_03102_),
    .A(net1053),
    .Y(_03103_));
 sg13g2_mux2_1 _09077_ (.A0(\dp.rf.rf[28][19] ),
    .A1(\dp.rf.rf[29][19] ),
    .S(net1321),
    .X(_03104_));
 sg13g2_nand3_1 _09078_ (.B(net1055),
    .C(_03104_),
    .A(net1067),
    .Y(_03105_));
 sg13g2_mux2_1 _09079_ (.A0(\dp.rf.rf[20][19] ),
    .A1(\dp.rf.rf[21][19] ),
    .S(net1326),
    .X(_03106_));
 sg13g2_nand3_1 _09080_ (.B(net1055),
    .C(_03106_),
    .A(net1060),
    .Y(_03107_));
 sg13g2_nand4_1 _09081_ (.B(_03103_),
    .C(_03105_),
    .A(_03101_),
    .Y(_03108_),
    .D(_03107_));
 sg13g2_nor4_2 _09082_ (.A(_03085_),
    .B(_03094_),
    .C(_03099_),
    .Y(_03109_),
    .D(_03108_));
 sg13g2_and2_1 _09083_ (.A(_03080_),
    .B(_03109_),
    .X(_03110_));
 sg13g2_buf_1 fanout1015 (.A(net1024),
    .X(net1015));
 sg13g2_nor2_1 _09085_ (.A(_02976_),
    .B(_03110_),
    .Y(net143));
 sg13g2_mux2_1 _09086_ (.A0(\dp.rf.rf[28][20] ),
    .A1(\dp.rf.rf[29][20] ),
    .S(net1324),
    .X(_03112_));
 sg13g2_nand3_1 _09087_ (.B(net1054),
    .C(_03112_),
    .A(net1067),
    .Y(_03113_));
 sg13g2_mux2_1 _09088_ (.A0(\dp.rf.rf[30][20] ),
    .A1(\dp.rf.rf[31][20] ),
    .S(net1340),
    .X(_03114_));
 sg13g2_nand2_1 _09089_ (.Y(_03115_),
    .A(_02663_),
    .B(_03114_));
 sg13g2_mux2_1 _09090_ (.A0(\dp.rf.rf[20][20] ),
    .A1(\dp.rf.rf[21][20] ),
    .S(net1335),
    .X(_03116_));
 sg13g2_nand3_1 _09091_ (.B(net1054),
    .C(_03116_),
    .A(net1060),
    .Y(_03117_));
 sg13g2_mux2_1 _09092_ (.A0(\dp.rf.rf[22][20] ),
    .A1(\dp.rf.rf[23][20] ),
    .S(net1311),
    .X(_03118_));
 sg13g2_nand3_1 _09093_ (.B(net1054),
    .C(_03118_),
    .A(net1053),
    .Y(_03119_));
 sg13g2_nand4_1 _09094_ (.B(_03115_),
    .C(_03117_),
    .A(_03113_),
    .Y(_03120_),
    .D(_03119_));
 sg13g2_buf_2 fanout1014 (.A(net1015),
    .X(net1014));
 sg13g2_mux4_1 _09096_ (.S0(net1335),
    .A0(\dp.rf.rf[24][20] ),
    .A1(\dp.rf.rf[25][20] ),
    .A2(\dp.rf.rf[26][20] ),
    .A3(\dp.rf.rf[27][20] ),
    .S1(net1286),
    .X(_03122_));
 sg13g2_nand2_1 _09097_ (.Y(_03123_),
    .A(net1265),
    .B(_03122_));
 sg13g2_mux4_1 _09098_ (.S0(net1335),
    .A0(\dp.rf.rf[16][20] ),
    .A1(\dp.rf.rf[17][20] ),
    .A2(\dp.rf.rf[18][20] ),
    .A3(\dp.rf.rf[19][20] ),
    .S1(net1286),
    .X(_03124_));
 sg13g2_nand2_1 _09099_ (.Y(_03125_),
    .A(net1046),
    .B(_03124_));
 sg13g2_buf_1 fanout1013 (.A(net1015),
    .X(net1013));
 sg13g2_inv_2 _09101_ (.Y(_03127_),
    .A(net1277));
 sg13g2_nand2_2 _09102_ (.Y(_03128_),
    .A(net1258),
    .B(_03127_));
 sg13g2_a21oi_1 _09103_ (.A1(_03123_),
    .A2(_03125_),
    .Y(_03129_),
    .B1(_03128_));
 sg13g2_buf_2 fanout1012 (.A(net1015),
    .X(net1012));
 sg13g2_buf_2 fanout1011 (.A(net1012),
    .X(net1011));
 sg13g2_buf_2 fanout1010 (.A(_03676_),
    .X(net1010));
 sg13g2_nor2b_1 _09107_ (.A(net1331),
    .B_N(\dp.rf.rf[10][20] ),
    .Y(_03133_));
 sg13g2_a22oi_1 _09108_ (.Y(_03134_),
    .B1(net1096),
    .B2(_03133_),
    .A2(\dp.rf.rf[11][20] ),
    .A1(net1331));
 sg13g2_buf_4 fanout1009 (.X(net1009),
    .A(net1010));
 sg13g2_nor2b_1 _09110_ (.A(net1332),
    .B_N(\dp.rf.rf[0][20] ),
    .Y(_03136_));
 sg13g2_a22oi_1 _09111_ (.Y(_03137_),
    .B1(net1081),
    .B2(_03136_),
    .A2(\dp.rf.rf[1][20] ),
    .A1(net1332));
 sg13g2_buf_4 fanout1008 (.X(net1008),
    .A(net1010));
 sg13g2_nor2b_1 _09113_ (.A(net1331),
    .B_N(\dp.rf.rf[8][20] ),
    .Y(_03139_));
 sg13g2_a22oi_1 _09114_ (.Y(_03140_),
    .B1(net1088),
    .B2(_03139_),
    .A2(\dp.rf.rf[9][20] ),
    .A1(net1331));
 sg13g2_buf_4 fanout1007 (.X(net1007),
    .A(net1008));
 sg13g2_mux2_1 _09116_ (.A0(\dp.rf.rf[2][20] ),
    .A1(\dp.rf.rf[3][20] ),
    .S(net1332),
    .X(_03142_));
 sg13g2_o21ai_1 _09117_ (.B1(net1050),
    .Y(_03143_),
    .A1(net1075),
    .A2(_03142_));
 sg13g2_nor4_1 _09118_ (.A(_03134_),
    .B(_03137_),
    .C(_03140_),
    .D(_03143_),
    .Y(_03144_));
 sg13g2_buf_4 fanout1006 (.X(net1006),
    .A(_03683_));
 sg13g2_nor2b_1 _09120_ (.A(net1332),
    .B_N(\dp.rf.rf[14][20] ),
    .Y(_03146_));
 sg13g2_a22oi_1 _09121_ (.Y(_03147_),
    .B1(net1100),
    .B2(_03146_),
    .A2(\dp.rf.rf[15][20] ),
    .A1(net1332));
 sg13g2_nor2b_1 _09122_ (.A(net1331),
    .B_N(\dp.rf.rf[6][20] ),
    .Y(_03148_));
 sg13g2_a22oi_1 _09123_ (.Y(_03149_),
    .B1(net1075),
    .B2(_03148_),
    .A2(\dp.rf.rf[7][20] ),
    .A1(net1331));
 sg13g2_nor2b_1 _09124_ (.A(net1333),
    .B_N(\dp.rf.rf[12][20] ),
    .Y(_03150_));
 sg13g2_a22oi_1 _09125_ (.Y(_03151_),
    .B1(net1088),
    .B2(_03150_),
    .A2(\dp.rf.rf[13][20] ),
    .A1(net1333));
 sg13g2_mux2_1 _09126_ (.A0(\dp.rf.rf[4][20] ),
    .A1(\dp.rf.rf[5][20] ),
    .S(net1331),
    .X(_03152_));
 sg13g2_o21ai_1 _09127_ (.B1(net1062),
    .Y(_03153_),
    .A1(net1081),
    .A2(_03152_));
 sg13g2_nor4_1 _09128_ (.A(_03147_),
    .B(_03149_),
    .C(_03151_),
    .D(_03153_),
    .Y(_03154_));
 sg13g2_nor4_2 _09129_ (.A(_03120_),
    .B(_03129_),
    .C(_03144_),
    .Y(_03155_),
    .D(_03154_));
 sg13g2_nor2_1 _09130_ (.A(_03050_),
    .B(_03155_),
    .Y(net145));
 sg13g2_mux4_1 _09131_ (.S0(net1310),
    .A0(\dp.rf.rf[12][21] ),
    .A1(\dp.rf.rf[13][21] ),
    .A2(\dp.rf.rf[14][21] ),
    .A3(\dp.rf.rf[15][21] ),
    .S1(net1280),
    .X(_03156_));
 sg13g2_mux4_1 _09132_ (.S0(net1310),
    .A0(\dp.rf.rf[4][21] ),
    .A1(\dp.rf.rf[5][21] ),
    .A2(\dp.rf.rf[6][21] ),
    .A3(\dp.rf.rf[7][21] ),
    .S1(net1280),
    .X(_03157_));
 sg13g2_and2_1 _09133_ (.A(net1044),
    .B(_03157_),
    .X(_03158_));
 sg13g2_a22oi_1 _09134_ (.Y(_03159_),
    .B1(_03158_),
    .B2(_02746_),
    .A2(_03156_),
    .A1(net1262));
 sg13g2_mux4_1 _09135_ (.S0(net1308),
    .A0(\dp.rf.rf[8][21] ),
    .A1(\dp.rf.rf[9][21] ),
    .A2(\dp.rf.rf[10][21] ),
    .A3(\dp.rf.rf[11][21] ),
    .S1(net1280),
    .X(_03160_));
 sg13g2_mux4_1 _09136_ (.S0(net1310),
    .A0(\dp.rf.rf[0][21] ),
    .A1(\dp.rf.rf[1][21] ),
    .A2(\dp.rf.rf[2][21] ),
    .A3(\dp.rf.rf[3][21] ),
    .S1(net1280),
    .X(_03161_));
 sg13g2_and2_1 _09137_ (.A(net1044),
    .B(_03161_),
    .X(_03162_));
 sg13g2_a22oi_1 _09138_ (.Y(_03163_),
    .B1(_03162_),
    .B2(net1105),
    .A2(_03160_),
    .A1(net1262));
 sg13g2_mux4_1 _09139_ (.S0(net1310),
    .A0(\dp.rf.rf[24][21] ),
    .A1(\dp.rf.rf[25][21] ),
    .A2(\dp.rf.rf[26][21] ),
    .A3(\dp.rf.rf[27][21] ),
    .S1(net1280),
    .X(_03164_));
 sg13g2_mux4_1 _09140_ (.S0(net1310),
    .A0(\dp.rf.rf[16][21] ),
    .A1(\dp.rf.rf[17][21] ),
    .A2(\dp.rf.rf[18][21] ),
    .A3(\dp.rf.rf[19][21] ),
    .S1(net1280),
    .X(_03165_));
 sg13g2_and2_1 _09141_ (.A(net1044),
    .B(_03165_),
    .X(_03166_));
 sg13g2_a22oi_1 _09142_ (.Y(_03167_),
    .B1(_03166_),
    .B2(_03128_),
    .A2(_03164_),
    .A1(net1263));
 sg13g2_mux2_1 _09143_ (.A0(\dp.rf.rf[22][21] ),
    .A1(\dp.rf.rf[23][21] ),
    .S(net1312),
    .X(_03168_));
 sg13g2_nor3_1 _09144_ (.A(net1073),
    .B(_02768_),
    .C(_03168_),
    .Y(_03169_));
 sg13g2_mux2_1 _09145_ (.A0(\dp.rf.rf[20][21] ),
    .A1(\dp.rf.rf[21][21] ),
    .S(net1312),
    .X(_03170_));
 sg13g2_nor3_1 _09146_ (.A(net1079),
    .B(_02768_),
    .C(_03170_),
    .Y(_03171_));
 sg13g2_nor2b_1 _09147_ (.A(net1312),
    .B_N(\dp.rf.rf[30][21] ),
    .Y(_03172_));
 sg13g2_a22oi_1 _09148_ (.Y(_03173_),
    .B1(_02822_),
    .B2(_03172_),
    .A2(\dp.rf.rf[31][21] ),
    .A1(net1312));
 sg13g2_mux2_1 _09149_ (.A0(\dp.rf.rf[28][21] ),
    .A1(\dp.rf.rf[29][21] ),
    .S(net1312),
    .X(_03174_));
 sg13g2_nor3_1 _09150_ (.A(net1086),
    .B(_02768_),
    .C(_03174_),
    .Y(_03175_));
 sg13g2_or4_1 _09151_ (.A(_03169_),
    .B(_03171_),
    .C(_03173_),
    .D(_03175_),
    .X(_03176_));
 sg13g2_nor4_2 _09152_ (.A(_03159_),
    .B(_03163_),
    .C(_03167_),
    .Y(_03177_),
    .D(_03176_));
 sg13g2_nor2b_1 _09153_ (.A(_03050_),
    .B_N(_03177_),
    .Y(net146));
 sg13g2_mux4_1 _09154_ (.S0(net1331),
    .A0(\dp.rf.rf[12][22] ),
    .A1(\dp.rf.rf[13][22] ),
    .A2(\dp.rf.rf[14][22] ),
    .A3(\dp.rf.rf[15][22] ),
    .S1(net1288),
    .X(_03178_));
 sg13g2_nand2_1 _09155_ (.Y(_03179_),
    .A(net1265),
    .B(_03178_));
 sg13g2_mux4_1 _09156_ (.S0(net1332),
    .A0(\dp.rf.rf[4][22] ),
    .A1(\dp.rf.rf[5][22] ),
    .A2(\dp.rf.rf[6][22] ),
    .A3(\dp.rf.rf[7][22] ),
    .S1(net1288),
    .X(_03180_));
 sg13g2_nand2_1 _09157_ (.Y(_03181_),
    .A(net1046),
    .B(_03180_));
 sg13g2_a21oi_1 _09158_ (.A1(_03179_),
    .A2(_03181_),
    .Y(_03182_),
    .B1(_02746_));
 sg13g2_mux4_1 _09159_ (.S0(net1334),
    .A0(\dp.rf.rf[20][22] ),
    .A1(\dp.rf.rf[21][22] ),
    .A2(\dp.rf.rf[22][22] ),
    .A3(\dp.rf.rf[23][22] ),
    .S1(net1286),
    .X(_03183_));
 sg13g2_mux4_1 _09160_ (.S0(net1335),
    .A0(\dp.rf.rf[28][22] ),
    .A1(\dp.rf.rf[29][22] ),
    .A2(\dp.rf.rf[30][22] ),
    .A3(\dp.rf.rf[31][22] ),
    .S1(net1287),
    .X(_03184_));
 sg13g2_nor2b_1 _09161_ (.A(net1042),
    .B_N(_03184_),
    .Y(_03185_));
 sg13g2_a21o_1 _09162_ (.A2(_03183_),
    .A1(net951),
    .B1(_03185_),
    .X(_03186_));
 sg13g2_buf_4 fanout1005 (.X(net1005),
    .A(_03689_));
 sg13g2_nor2b_1 _09164_ (.A(net1334),
    .B_N(\dp.rf.rf[26][22] ),
    .Y(_03188_));
 sg13g2_a22oi_1 _09165_ (.Y(_03189_),
    .B1(net1096),
    .B2(_03188_),
    .A2(\dp.rf.rf[27][22] ),
    .A1(net1334));
 sg13g2_nor2b_1 _09166_ (.A(net1334),
    .B_N(\dp.rf.rf[16][22] ),
    .Y(_03190_));
 sg13g2_a22oi_1 _09167_ (.Y(_03191_),
    .B1(net1081),
    .B2(_03190_),
    .A2(\dp.rf.rf[17][22] ),
    .A1(net1334));
 sg13g2_nor2b_1 _09168_ (.A(net1334),
    .B_N(\dp.rf.rf[24][22] ),
    .Y(_03192_));
 sg13g2_a22oi_1 _09169_ (.Y(_03193_),
    .B1(net1088),
    .B2(_03192_),
    .A2(\dp.rf.rf[25][22] ),
    .A1(net1334));
 sg13g2_mux2_1 _09170_ (.A0(\dp.rf.rf[18][22] ),
    .A1(\dp.rf.rf[19][22] ),
    .S(net1334),
    .X(_03194_));
 sg13g2_o21ai_1 _09171_ (.B1(net1072),
    .Y(_03195_),
    .A1(net1075),
    .A2(_03194_));
 sg13g2_nor4_1 _09172_ (.A(_03189_),
    .B(_03191_),
    .C(_03193_),
    .D(_03195_),
    .Y(_03196_));
 sg13g2_nor2b_1 _09173_ (.A(net1336),
    .B_N(\dp.rf.rf[2][22] ),
    .Y(_03197_));
 sg13g2_a22oi_1 _09174_ (.Y(_03198_),
    .B1(net1075),
    .B2(_03197_),
    .A2(\dp.rf.rf[3][22] ),
    .A1(net1336));
 sg13g2_nor2b_1 _09175_ (.A(net1336),
    .B_N(\dp.rf.rf[0][22] ),
    .Y(_03199_));
 sg13g2_a22oi_1 _09176_ (.Y(_03200_),
    .B1(net1081),
    .B2(_03199_),
    .A2(\dp.rf.rf[1][22] ),
    .A1(net1337));
 sg13g2_nor2b_1 _09177_ (.A(net1336),
    .B_N(\dp.rf.rf[10][22] ),
    .Y(_03201_));
 sg13g2_a22oi_1 _09178_ (.Y(_03202_),
    .B1(net1096),
    .B2(_03201_),
    .A2(\dp.rf.rf[11][22] ),
    .A1(net1336));
 sg13g2_mux2_1 _09179_ (.A0(\dp.rf.rf[8][22] ),
    .A1(\dp.rf.rf[9][22] ),
    .S(net1336),
    .X(_03203_));
 sg13g2_o21ai_1 _09180_ (.B1(net1050),
    .Y(_03204_),
    .A1(net1088),
    .A2(_03203_));
 sg13g2_nor4_1 _09181_ (.A(_03198_),
    .B(_03200_),
    .C(_03202_),
    .D(_03204_),
    .Y(_03205_));
 sg13g2_nor4_2 _09182_ (.A(_03182_),
    .B(_03186_),
    .C(_03196_),
    .Y(_03206_),
    .D(_03205_));
 sg13g2_nor2_1 _09183_ (.A(_03050_),
    .B(_03206_),
    .Y(net147));
 sg13g2_mux4_1 _09184_ (.S0(net1315),
    .A0(\dp.rf.rf[20][23] ),
    .A1(\dp.rf.rf[21][23] ),
    .A2(\dp.rf.rf[22][23] ),
    .A3(\dp.rf.rf[23][23] ),
    .S1(net1282),
    .X(_03207_));
 sg13g2_mux4_1 _09185_ (.S0(net1315),
    .A0(\dp.rf.rf[28][23] ),
    .A1(\dp.rf.rf[29][23] ),
    .A2(\dp.rf.rf[30][23] ),
    .A3(\dp.rf.rf[31][23] ),
    .S1(net1282),
    .X(_03208_));
 sg13g2_nor2b_1 _09186_ (.A(net1042),
    .B_N(_03208_),
    .Y(_03209_));
 sg13g2_a21o_1 _09187_ (.A2(_03207_),
    .A1(net951),
    .B1(_03209_),
    .X(_03210_));
 sg13g2_mux4_1 _09188_ (.S0(net1325),
    .A0(\dp.rf.rf[2][23] ),
    .A1(\dp.rf.rf[3][23] ),
    .A2(\dp.rf.rf[10][23] ),
    .A3(\dp.rf.rf[11][23] ),
    .S1(net1264),
    .X(_03211_));
 sg13g2_nand2_1 _09189_ (.Y(_03212_),
    .A(net1284),
    .B(_03211_));
 sg13g2_mux4_1 _09190_ (.S0(net1325),
    .A0(\dp.rf.rf[0][23] ),
    .A1(\dp.rf.rf[1][23] ),
    .A2(\dp.rf.rf[8][23] ),
    .A3(\dp.rf.rf[9][23] ),
    .S1(net1264),
    .X(_03213_));
 sg13g2_nand2_1 _09191_ (.Y(_03214_),
    .A(net1101),
    .B(_03213_));
 sg13g2_nand2b_1 _09192_ (.Y(_03215_),
    .B(net1051),
    .A_N(_02592_));
 sg13g2_a21oi_1 _09193_ (.A1(_03212_),
    .A2(_03214_),
    .Y(_03216_),
    .B1(_03215_));
 sg13g2_nor2b_1 _09194_ (.A(net1316),
    .B_N(\dp.rf.rf[14][23] ),
    .Y(_03217_));
 sg13g2_a22oi_1 _09195_ (.Y(_03218_),
    .B1(net1095),
    .B2(_03217_),
    .A2(\dp.rf.rf[15][23] ),
    .A1(net1316));
 sg13g2_buf_4 fanout1004 (.X(net1004),
    .A(net1005));
 sg13g2_nor2b_1 _09197_ (.A(net1316),
    .B_N(\dp.rf.rf[12][23] ),
    .Y(_03220_));
 sg13g2_a22oi_1 _09198_ (.Y(_03221_),
    .B1(net1087),
    .B2(_03220_),
    .A2(\dp.rf.rf[13][23] ),
    .A1(net1316));
 sg13g2_nor2b_1 _09199_ (.A(net1316),
    .B_N(\dp.rf.rf[4][23] ),
    .Y(_03222_));
 sg13g2_a22oi_1 _09200_ (.Y(_03223_),
    .B1(net1080),
    .B2(_03222_),
    .A2(\dp.rf.rf[5][23] ),
    .A1(net1316));
 sg13g2_mux2_1 _09201_ (.A0(\dp.rf.rf[6][23] ),
    .A1(\dp.rf.rf[7][23] ),
    .S(net1318),
    .X(_03224_));
 sg13g2_o21ai_1 _09202_ (.B1(net1061),
    .Y(_03225_),
    .A1(net1074),
    .A2(_03224_));
 sg13g2_nor4_1 _09203_ (.A(_03218_),
    .B(_03221_),
    .C(_03223_),
    .D(_03225_),
    .Y(_03226_));
 sg13g2_nor2b_1 _09204_ (.A(net1317),
    .B_N(\dp.rf.rf[18][23] ),
    .Y(_03227_));
 sg13g2_a22oi_1 _09205_ (.Y(_03228_),
    .B1(net1073),
    .B2(_03227_),
    .A2(\dp.rf.rf[19][23] ),
    .A1(net1317));
 sg13g2_nor2b_1 _09206_ (.A(net1317),
    .B_N(\dp.rf.rf[16][23] ),
    .Y(_03229_));
 sg13g2_a22oi_1 _09207_ (.Y(_03230_),
    .B1(net1080),
    .B2(_03229_),
    .A2(\dp.rf.rf[17][23] ),
    .A1(net1317));
 sg13g2_nor2b_1 _09208_ (.A(net1317),
    .B_N(\dp.rf.rf[26][23] ),
    .Y(_03231_));
 sg13g2_a22oi_1 _09209_ (.Y(_03232_),
    .B1(net1096),
    .B2(_03231_),
    .A2(\dp.rf.rf[27][23] ),
    .A1(net1317));
 sg13g2_mux2_1 _09210_ (.A0(\dp.rf.rf[24][23] ),
    .A1(\dp.rf.rf[25][23] ),
    .S(net1317),
    .X(_03233_));
 sg13g2_o21ai_1 _09211_ (.B1(net1069),
    .Y(_03234_),
    .A1(net1087),
    .A2(_03233_));
 sg13g2_nor4_1 _09212_ (.A(_03228_),
    .B(_03230_),
    .C(_03232_),
    .D(_03234_),
    .Y(_03235_));
 sg13g2_nor4_2 _09213_ (.A(_03210_),
    .B(_03216_),
    .C(_03226_),
    .Y(_03236_),
    .D(_03235_));
 sg13g2_nor2_1 _09214_ (.A(net913),
    .B(_03236_),
    .Y(net148));
 sg13g2_buf_4 fanout1003 (.X(net1003),
    .A(_03715_));
 sg13g2_nor2b_1 _09216_ (.A(net1308),
    .B_N(\dp.rf.rf[6][24] ),
    .Y(_03238_));
 sg13g2_a22oi_1 _09217_ (.Y(_03239_),
    .B1(net1073),
    .B2(_03238_),
    .A2(\dp.rf.rf[7][24] ),
    .A1(net1308));
 sg13g2_nor2b_1 _09218_ (.A(net1308),
    .B_N(\dp.rf.rf[4][24] ),
    .Y(_03240_));
 sg13g2_a22oi_1 _09219_ (.Y(_03241_),
    .B1(net1079),
    .B2(_03240_),
    .A2(\dp.rf.rf[5][24] ),
    .A1(net1308));
 sg13g2_nor2b_1 _09220_ (.A(net1308),
    .B_N(\dp.rf.rf[14][24] ),
    .Y(_03242_));
 sg13g2_a22oi_1 _09221_ (.Y(_03243_),
    .B1(net1096),
    .B2(_03242_),
    .A2(\dp.rf.rf[15][24] ),
    .A1(net1308));
 sg13g2_mux2_1 _09222_ (.A0(\dp.rf.rf[12][24] ),
    .A1(\dp.rf.rf[13][24] ),
    .S(net1308),
    .X(_03244_));
 sg13g2_o21ai_1 _09223_ (.B1(net1061),
    .Y(_03245_),
    .A1(net1088),
    .A2(_03244_));
 sg13g2_or4_1 _09224_ (.A(_03239_),
    .B(_03241_),
    .C(_03243_),
    .D(_03245_),
    .X(_03246_));
 sg13g2_mux4_1 _09225_ (.S0(net1309),
    .A0(\dp.rf.rf[18][24] ),
    .A1(\dp.rf.rf[19][24] ),
    .A2(\dp.rf.rf[26][24] ),
    .A3(\dp.rf.rf[27][24] ),
    .S1(net1263),
    .X(_03247_));
 sg13g2_nor2_1 _09226_ (.A(net1101),
    .B(_03247_),
    .Y(_03248_));
 sg13g2_nor2b_1 _09227_ (.A(net1311),
    .B_N(\dp.rf.rf[24][24] ),
    .Y(_03249_));
 sg13g2_a22oi_1 _09228_ (.Y(_03250_),
    .B1(net1088),
    .B2(_03249_),
    .A2(\dp.rf.rf[25][24] ),
    .A1(net1309));
 sg13g2_buf_2 fanout1002 (.A(net1003),
    .X(net1002));
 sg13g2_nor2b_1 _09230_ (.A(net1309),
    .B_N(\dp.rf.rf[16][24] ),
    .Y(_03252_));
 sg13g2_a22oi_1 _09231_ (.Y(_03253_),
    .B1(net1079),
    .B2(_03252_),
    .A2(\dp.rf.rf[17][24] ),
    .A1(net1309));
 sg13g2_or4_1 _09232_ (.A(_03128_),
    .B(_03248_),
    .C(_03250_),
    .D(_03253_),
    .X(_03254_));
 sg13g2_mux2_1 _09233_ (.A0(\dp.rf.rf[10][24] ),
    .A1(\dp.rf.rf[11][24] ),
    .S(net1330),
    .X(_03255_));
 sg13g2_mux2_1 _09234_ (.A0(\dp.rf.rf[2][24] ),
    .A1(\dp.rf.rf[3][24] ),
    .S(net1330),
    .X(_03256_));
 sg13g2_mux2_1 _09235_ (.A0(\dp.rf.rf[8][24] ),
    .A1(\dp.rf.rf[9][24] ),
    .S(net1330),
    .X(_03257_));
 sg13g2_and2_1 _09236_ (.A(net1330),
    .B(\dp.rf.rf[1][24] ),
    .X(_03258_));
 sg13g2_mux4_1 _09237_ (.S0(net1046),
    .A0(_03255_),
    .A1(_03256_),
    .A2(_03257_),
    .A3(_03258_),
    .S1(net1101),
    .X(_03259_));
 sg13g2_mux4_1 _09238_ (.S0(net1330),
    .A0(\dp.rf.rf[20][24] ),
    .A1(\dp.rf.rf[21][24] ),
    .A2(\dp.rf.rf[22][24] ),
    .A3(\dp.rf.rf[23][24] ),
    .S1(net1286),
    .X(_03260_));
 sg13g2_mux4_1 _09239_ (.S0(net1311),
    .A0(\dp.rf.rf[28][24] ),
    .A1(\dp.rf.rf[29][24] ),
    .A2(\dp.rf.rf[30][24] ),
    .A3(\dp.rf.rf[31][24] ),
    .S1(net1280),
    .X(_03261_));
 sg13g2_nor2b_1 _09240_ (.A(net1042),
    .B_N(_03261_),
    .Y(_03262_));
 sg13g2_a221oi_1 _09241_ (.B2(net951),
    .C1(_03262_),
    .B1(_03260_),
    .A1(net1050),
    .Y(_03263_),
    .A2(_03259_));
 sg13g2_and3_1 _09242_ (.X(_03264_),
    .A(_03246_),
    .B(_03254_),
    .C(_03263_));
 sg13g2_buf_4 fanout1001 (.X(net1001),
    .A(_03725_));
 sg13g2_nor2_1 _09244_ (.A(net913),
    .B(_03264_),
    .Y(net149));
 sg13g2_buf_2 fanout1000 (.A(net1001),
    .X(net1000));
 sg13g2_mux4_1 _09246_ (.S0(net1305),
    .A0(\dp.rf.rf[20][25] ),
    .A1(\dp.rf.rf[21][25] ),
    .A2(\dp.rf.rf[22][25] ),
    .A3(\dp.rf.rf[23][25] ),
    .S1(net1279),
    .X(_03267_));
 sg13g2_mux4_1 _09247_ (.S0(net1306),
    .A0(\dp.rf.rf[28][25] ),
    .A1(\dp.rf.rf[29][25] ),
    .A2(\dp.rf.rf[30][25] ),
    .A3(\dp.rf.rf[31][25] ),
    .S1(net1278),
    .X(_03268_));
 sg13g2_nor2b_1 _09248_ (.A(net1042),
    .B_N(_03268_),
    .Y(_03269_));
 sg13g2_a21o_1 _09249_ (.A2(_03267_),
    .A1(net951),
    .B1(_03269_),
    .X(_03270_));
 sg13g2_nor2b_1 _09250_ (.A(net1305),
    .B_N(\dp.rf.rf[6][25] ),
    .Y(_03271_));
 sg13g2_a22oi_1 _09251_ (.Y(_03272_),
    .B1(net1073),
    .B2(_03271_),
    .A2(\dp.rf.rf[7][25] ),
    .A1(net1305));
 sg13g2_nor2b_1 _09252_ (.A(net1303),
    .B_N(\dp.rf.rf[14][25] ),
    .Y(_03273_));
 sg13g2_a22oi_1 _09253_ (.Y(_03274_),
    .B1(net1095),
    .B2(_03273_),
    .A2(\dp.rf.rf[15][25] ),
    .A1(net1303));
 sg13g2_nor2b_1 _09254_ (.A(net1305),
    .B_N(\dp.rf.rf[4][25] ),
    .Y(_03275_));
 sg13g2_a22oi_1 _09255_ (.Y(_03276_),
    .B1(net1079),
    .B2(_03275_),
    .A2(\dp.rf.rf[5][25] ),
    .A1(net1305));
 sg13g2_mux2_1 _09256_ (.A0(\dp.rf.rf[12][25] ),
    .A1(\dp.rf.rf[13][25] ),
    .S(net1303),
    .X(_03277_));
 sg13g2_o21ai_1 _09257_ (.B1(net1061),
    .Y(_03278_),
    .A1(net1086),
    .A2(_03277_));
 sg13g2_nor4_1 _09258_ (.A(_03272_),
    .B(_03274_),
    .C(_03276_),
    .D(_03278_),
    .Y(_03279_));
 sg13g2_nor2b_1 _09259_ (.A(net1305),
    .B_N(\dp.rf.rf[18][25] ),
    .Y(_03280_));
 sg13g2_a22oi_1 _09260_ (.Y(_03281_),
    .B1(net1073),
    .B2(_03280_),
    .A2(\dp.rf.rf[19][25] ),
    .A1(net1303));
 sg13g2_buf_1 fanout999 (.A(net1000),
    .X(net999));
 sg13g2_nor2b_1 _09262_ (.A(net1303),
    .B_N(\dp.rf.rf[26][25] ),
    .Y(_03283_));
 sg13g2_a22oi_1 _09263_ (.Y(_03284_),
    .B1(net1095),
    .B2(_03283_),
    .A2(\dp.rf.rf[27][25] ),
    .A1(net1303));
 sg13g2_nor2b_1 _09264_ (.A(net1304),
    .B_N(\dp.rf.rf[16][25] ),
    .Y(_03285_));
 sg13g2_a22oi_1 _09265_ (.Y(_03286_),
    .B1(net1079),
    .B2(_03285_),
    .A2(\dp.rf.rf[17][25] ),
    .A1(net1304));
 sg13g2_mux2_1 _09266_ (.A0(\dp.rf.rf[24][25] ),
    .A1(\dp.rf.rf[25][25] ),
    .S(net1307),
    .X(_03287_));
 sg13g2_o21ai_1 _09267_ (.B1(net1069),
    .Y(_03288_),
    .A1(net1086),
    .A2(_03287_));
 sg13g2_nor4_1 _09268_ (.A(_03281_),
    .B(_03284_),
    .C(_03286_),
    .D(_03288_),
    .Y(_03289_));
 sg13g2_mux4_1 _09269_ (.S0(net1303),
    .A0(\dp.rf.rf[2][25] ),
    .A1(\dp.rf.rf[3][25] ),
    .A2(\dp.rf.rf[10][25] ),
    .A3(\dp.rf.rf[11][25] ),
    .S1(net1262),
    .X(_03290_));
 sg13g2_nor2_1 _09270_ (.A(net1101),
    .B(_03290_),
    .Y(_03291_));
 sg13g2_mux2_1 _09271_ (.A0(\dp.rf.rf[1][25] ),
    .A1(\dp.rf.rf[9][25] ),
    .S(net1262),
    .X(_03292_));
 sg13g2_buf_2 fanout998 (.A(net1000),
    .X(net998));
 sg13g2_a221oi_1 _09273_ (.B2(net1303),
    .C1(net1279),
    .B1(_03292_),
    .A1(\dp.rf.rf[8][25] ),
    .Y(_03294_),
    .A2(_02731_));
 sg13g2_nor3_1 _09274_ (.A(net1105),
    .B(_03291_),
    .C(_03294_),
    .Y(_03295_));
 sg13g2_nor4_2 _09275_ (.A(_03270_),
    .B(_03279_),
    .C(_03289_),
    .Y(_03296_),
    .D(_03295_));
 sg13g2_nor2_1 _09276_ (.A(net913),
    .B(_03296_),
    .Y(net150));
 sg13g2_buf_2 fanout997 (.A(_03734_),
    .X(net997));
 sg13g2_mux4_1 _09278_ (.S0(net1330),
    .A0(\dp.rf.rf[8][26] ),
    .A1(\dp.rf.rf[9][26] ),
    .A2(\dp.rf.rf[10][26] ),
    .A3(\dp.rf.rf[11][26] ),
    .S1(net1286),
    .X(_03298_));
 sg13g2_mux4_1 _09279_ (.S0(net1330),
    .A0(\dp.rf.rf[0][26] ),
    .A1(\dp.rf.rf[1][26] ),
    .A2(\dp.rf.rf[2][26] ),
    .A3(\dp.rf.rf[3][26] ),
    .S1(net1286),
    .X(_03299_));
 sg13g2_mux4_1 _09280_ (.S0(net1330),
    .A0(\dp.rf.rf[12][26] ),
    .A1(\dp.rf.rf[13][26] ),
    .A2(\dp.rf.rf[14][26] ),
    .A3(\dp.rf.rf[15][26] ),
    .S1(net1286),
    .X(_03300_));
 sg13g2_mux4_1 _09281_ (.S0(net1333),
    .A0(\dp.rf.rf[4][26] ),
    .A1(\dp.rf.rf[5][26] ),
    .A2(\dp.rf.rf[6][26] ),
    .A3(\dp.rf.rf[7][26] ),
    .S1(net1286),
    .X(_03301_));
 sg13g2_buf_1 fanout996 (.A(net997),
    .X(net996));
 sg13g2_mux4_1 _09283_ (.S0(net1046),
    .A0(_03298_),
    .A1(_03299_),
    .A2(_03300_),
    .A3(_03301_),
    .S1(net1275),
    .X(_03303_));
 sg13g2_and2_1 _09284_ (.A(net1051),
    .B(_02592_),
    .X(_03304_));
 sg13g2_buf_4 fanout995 (.X(net995),
    .A(net997));
 sg13g2_buf_2 fanout994 (.A(_03745_),
    .X(net994));
 sg13g2_nor2_1 _09287_ (.A(net1259),
    .B(net949),
    .Y(_03307_));
 sg13g2_mux4_1 _09288_ (.S0(net1306),
    .A0(\dp.rf.rf[24][26] ),
    .A1(\dp.rf.rf[25][26] ),
    .A2(\dp.rf.rf[26][26] ),
    .A3(\dp.rf.rf[27][26] ),
    .S1(net1278),
    .X(_03308_));
 sg13g2_mux4_1 _09289_ (.S0(net1306),
    .A0(\dp.rf.rf[16][26] ),
    .A1(\dp.rf.rf[17][26] ),
    .A2(\dp.rf.rf[18][26] ),
    .A3(\dp.rf.rf[19][26] ),
    .S1(net1278),
    .X(_03309_));
 sg13g2_mux4_1 _09290_ (.S0(net1306),
    .A0(\dp.rf.rf[28][26] ),
    .A1(\dp.rf.rf[29][26] ),
    .A2(\dp.rf.rf[30][26] ),
    .A3(\dp.rf.rf[31][26] ),
    .S1(net1278),
    .X(_03310_));
 sg13g2_mux4_1 _09291_ (.S0(net1306),
    .A0(\dp.rf.rf[20][26] ),
    .A1(\dp.rf.rf[21][26] ),
    .A2(\dp.rf.rf[22][26] ),
    .A3(\dp.rf.rf[23][26] ),
    .S1(net1278),
    .X(_03311_));
 sg13g2_mux4_1 _09292_ (.S0(net1044),
    .A0(_03308_),
    .A1(_03309_),
    .A2(_03310_),
    .A3(_03311_),
    .S1(net15),
    .X(_03312_));
 sg13g2_and2_1 _09293_ (.A(net1259),
    .B(_03312_),
    .X(_03313_));
 sg13g2_a21oi_2 _09294_ (.B1(_03313_),
    .Y(_03314_),
    .A2(_03307_),
    .A1(_03303_));
 sg13g2_nor2_1 _09295_ (.A(net913),
    .B(_03314_),
    .Y(net151));
 sg13g2_mux4_1 _09296_ (.S0(net1312),
    .A0(\dp.rf.rf[12][27] ),
    .A1(\dp.rf.rf[13][27] ),
    .A2(\dp.rf.rf[14][27] ),
    .A3(\dp.rf.rf[15][27] ),
    .S1(net1280),
    .X(_03315_));
 sg13g2_mux4_1 _09297_ (.S0(net1325),
    .A0(\dp.rf.rf[4][27] ),
    .A1(\dp.rf.rf[5][27] ),
    .A2(\dp.rf.rf[6][27] ),
    .A3(\dp.rf.rf[7][27] ),
    .S1(net1284),
    .X(_03316_));
 sg13g2_and2_1 _09298_ (.A(net1044),
    .B(_03316_),
    .X(_03317_));
 sg13g2_a22oi_1 _09299_ (.Y(_03318_),
    .B1(_03317_),
    .B2(_02746_),
    .A2(_03315_),
    .A1(net1263));
 sg13g2_mux4_1 _09300_ (.S0(net1306),
    .A0(\dp.rf.rf[24][27] ),
    .A1(\dp.rf.rf[25][27] ),
    .A2(\dp.rf.rf[26][27] ),
    .A3(\dp.rf.rf[27][27] ),
    .S1(net1282),
    .X(_03319_));
 sg13g2_mux4_1 _09301_ (.S0(net1307),
    .A0(\dp.rf.rf[16][27] ),
    .A1(\dp.rf.rf[17][27] ),
    .A2(\dp.rf.rf[18][27] ),
    .A3(\dp.rf.rf[19][27] ),
    .S1(net1278),
    .X(_03320_));
 sg13g2_and2_1 _09302_ (.A(net1044),
    .B(_03320_),
    .X(_03321_));
 sg13g2_a22oi_1 _09303_ (.Y(_03322_),
    .B1(_03321_),
    .B2(_03128_),
    .A2(_03319_),
    .A1(net1262));
 sg13g2_mux4_1 _09304_ (.S0(net1306),
    .A0(\dp.rf.rf[28][27] ),
    .A1(\dp.rf.rf[29][27] ),
    .A2(\dp.rf.rf[30][27] ),
    .A3(\dp.rf.rf[31][27] ),
    .S1(net1278),
    .X(_03323_));
 sg13g2_mux4_1 _09305_ (.S0(net1306),
    .A0(\dp.rf.rf[20][27] ),
    .A1(\dp.rf.rf[21][27] ),
    .A2(\dp.rf.rf[22][27] ),
    .A3(\dp.rf.rf[23][27] ),
    .S1(net1282),
    .X(_03324_));
 sg13g2_and2_1 _09306_ (.A(net1044),
    .B(_03324_),
    .X(_03325_));
 sg13g2_a22oi_1 _09307_ (.Y(_03326_),
    .B1(_03325_),
    .B2(_02768_),
    .A2(_03323_),
    .A1(net1262));
 sg13g2_mux4_1 _09308_ (.S0(net1307),
    .A0(\dp.rf.rf[8][27] ),
    .A1(\dp.rf.rf[9][27] ),
    .A2(\dp.rf.rf[10][27] ),
    .A3(\dp.rf.rf[11][27] ),
    .S1(net1278),
    .X(_03327_));
 sg13g2_mux4_1 _09309_ (.S0(net1325),
    .A0(\dp.rf.rf[0][27] ),
    .A1(\dp.rf.rf[1][27] ),
    .A2(\dp.rf.rf[2][27] ),
    .A3(\dp.rf.rf[3][27] ),
    .S1(net1284),
    .X(_03328_));
 sg13g2_and2_1 _09310_ (.A(net1044),
    .B(_03328_),
    .X(_03329_));
 sg13g2_a22oi_1 _09311_ (.Y(_03330_),
    .B1(_03329_),
    .B2(net1105),
    .A2(_03327_),
    .A1(net1262));
 sg13g2_nor4_2 _09312_ (.A(_03318_),
    .B(_03322_),
    .C(_03326_),
    .Y(_03331_),
    .D(_03330_));
 sg13g2_nor2b_1 _09313_ (.A(_03050_),
    .B_N(_03331_),
    .Y(net152));
 sg13g2_mux4_1 _09314_ (.S0(net1312),
    .A0(\dp.rf.rf[20][28] ),
    .A1(\dp.rf.rf[21][28] ),
    .A2(\dp.rf.rf[22][28] ),
    .A3(\dp.rf.rf[23][28] ),
    .S1(net1281),
    .X(_03332_));
 sg13g2_mux4_1 _09315_ (.S0(net1307),
    .A0(\dp.rf.rf[28][28] ),
    .A1(\dp.rf.rf[29][28] ),
    .A2(\dp.rf.rf[30][28] ),
    .A3(\dp.rf.rf[31][28] ),
    .S1(net1279),
    .X(_03333_));
 sg13g2_nor2b_1 _09316_ (.A(net1042),
    .B_N(_03333_),
    .Y(_03334_));
 sg13g2_a21o_1 _09317_ (.A2(_03332_),
    .A1(net951),
    .B1(_03334_),
    .X(_03335_));
 sg13g2_mux4_1 _09318_ (.S0(net1311),
    .A0(\dp.rf.rf[2][28] ),
    .A1(\dp.rf.rf[3][28] ),
    .A2(\dp.rf.rf[10][28] ),
    .A3(\dp.rf.rf[11][28] ),
    .S1(net1263),
    .X(_03336_));
 sg13g2_nand2_1 _09319_ (.Y(_03337_),
    .A(net1281),
    .B(_03336_));
 sg13g2_mux4_1 _09320_ (.S0(net1313),
    .A0(\dp.rf.rf[0][28] ),
    .A1(\dp.rf.rf[1][28] ),
    .A2(\dp.rf.rf[8][28] ),
    .A3(\dp.rf.rf[9][28] ),
    .S1(net1263),
    .X(_03338_));
 sg13g2_nand2_1 _09321_ (.Y(_03339_),
    .A(net1101),
    .B(_03338_));
 sg13g2_a21oi_1 _09322_ (.A1(_03337_),
    .A2(_03339_),
    .Y(_03340_),
    .B1(_03215_));
 sg13g2_nor2b_1 _09323_ (.A(net1307),
    .B_N(\dp.rf.rf[6][28] ),
    .Y(_03341_));
 sg13g2_a22oi_1 _09324_ (.Y(_03342_),
    .B1(net1073),
    .B2(_03341_),
    .A2(\dp.rf.rf[7][28] ),
    .A1(net1307));
 sg13g2_nor2b_1 _09325_ (.A(net1307),
    .B_N(\dp.rf.rf[4][28] ),
    .Y(_03343_));
 sg13g2_a22oi_1 _09326_ (.Y(_03344_),
    .B1(net1079),
    .B2(_03343_),
    .A2(\dp.rf.rf[5][28] ),
    .A1(net1307));
 sg13g2_nor2b_1 _09327_ (.A(net1304),
    .B_N(\dp.rf.rf[14][28] ),
    .Y(_03345_));
 sg13g2_a22oi_1 _09328_ (.Y(_03346_),
    .B1(net1095),
    .B2(_03345_),
    .A2(\dp.rf.rf[15][28] ),
    .A1(net1304));
 sg13g2_mux2_1 _09329_ (.A0(\dp.rf.rf[12][28] ),
    .A1(\dp.rf.rf[13][28] ),
    .S(net1304),
    .X(_03347_));
 sg13g2_o21ai_1 _09330_ (.B1(net1061),
    .Y(_03348_),
    .A1(net1086),
    .A2(_03347_));
 sg13g2_nor4_1 _09331_ (.A(_03342_),
    .B(_03344_),
    .C(_03346_),
    .D(_03348_),
    .Y(_03349_));
 sg13g2_nor2b_1 _09332_ (.A(net1311),
    .B_N(\dp.rf.rf[18][28] ),
    .Y(_03350_));
 sg13g2_a22oi_1 _09333_ (.Y(_03351_),
    .B1(net1073),
    .B2(_03350_),
    .A2(\dp.rf.rf[19][28] ),
    .A1(net1311));
 sg13g2_nor2b_1 _09334_ (.A(net1311),
    .B_N(\dp.rf.rf[16][28] ),
    .Y(_03352_));
 sg13g2_a22oi_1 _09335_ (.Y(_03353_),
    .B1(net1079),
    .B2(_03352_),
    .A2(\dp.rf.rf[17][28] ),
    .A1(net1311));
 sg13g2_nor2b_1 _09336_ (.A(net1310),
    .B_N(\dp.rf.rf[26][28] ),
    .Y(_03354_));
 sg13g2_a22oi_1 _09337_ (.Y(_03355_),
    .B1(net1095),
    .B2(_03354_),
    .A2(\dp.rf.rf[27][28] ),
    .A1(net1309));
 sg13g2_mux2_1 _09338_ (.A0(\dp.rf.rf[24][28] ),
    .A1(\dp.rf.rf[25][28] ),
    .S(net1312),
    .X(_03356_));
 sg13g2_o21ai_1 _09339_ (.B1(net1069),
    .Y(_03357_),
    .A1(net1086),
    .A2(_03356_));
 sg13g2_nor4_1 _09340_ (.A(_03351_),
    .B(_03353_),
    .C(_03355_),
    .D(_03357_),
    .Y(_03358_));
 sg13g2_nor4_2 _09341_ (.A(_03335_),
    .B(_03340_),
    .C(_03349_),
    .Y(_03359_),
    .D(_03358_));
 sg13g2_nor2_1 _09342_ (.A(net913),
    .B(_03359_),
    .Y(net153));
 sg13g2_mux2_1 _09343_ (.A0(\dp.rf.rf[8][29] ),
    .A1(\dp.rf.rf[9][29] ),
    .S(net1337),
    .X(_03360_));
 sg13g2_mux2_1 _09344_ (.A0(\dp.rf.rf[10][29] ),
    .A1(\dp.rf.rf[11][29] ),
    .S(net1337),
    .X(_03361_));
 sg13g2_and2_1 _09345_ (.A(net1337),
    .B(\dp.rf.rf[1][29] ),
    .X(_03362_));
 sg13g2_mux2_1 _09346_ (.A0(\dp.rf.rf[2][29] ),
    .A1(\dp.rf.rf[3][29] ),
    .S(net1336),
    .X(_03363_));
 sg13g2_mux4_1 _09347_ (.S0(net1288),
    .A0(_03360_),
    .A1(_03361_),
    .A2(_03362_),
    .A3(_03363_),
    .S1(net1047),
    .X(_03364_));
 sg13g2_mux4_1 _09348_ (.S0(net1336),
    .A0(\dp.rf.rf[12][29] ),
    .A1(\dp.rf.rf[13][29] ),
    .A2(\dp.rf.rf[14][29] ),
    .A3(\dp.rf.rf[15][29] ),
    .S1(net1288),
    .X(_03365_));
 sg13g2_nand2_1 _09349_ (.Y(_03366_),
    .A(net1265),
    .B(_03365_));
 sg13g2_mux4_1 _09350_ (.S0(net1337),
    .A0(\dp.rf.rf[4][29] ),
    .A1(\dp.rf.rf[5][29] ),
    .A2(\dp.rf.rf[6][29] ),
    .A3(\dp.rf.rf[7][29] ),
    .S1(net1288),
    .X(_03367_));
 sg13g2_nand2_1 _09351_ (.Y(_03368_),
    .A(net1046),
    .B(_03367_));
 sg13g2_a21oi_1 _09352_ (.A1(_03366_),
    .A2(_03368_),
    .Y(_03369_),
    .B1(_02746_));
 sg13g2_mux4_1 _09353_ (.S0(net1335),
    .A0(\dp.rf.rf[24][29] ),
    .A1(\dp.rf.rf[25][29] ),
    .A2(\dp.rf.rf[26][29] ),
    .A3(\dp.rf.rf[27][29] ),
    .S1(net1287),
    .X(_03370_));
 sg13g2_mux4_1 _09354_ (.S0(net1335),
    .A0(\dp.rf.rf[16][29] ),
    .A1(\dp.rf.rf[17][29] ),
    .A2(\dp.rf.rf[18][29] ),
    .A3(\dp.rf.rf[19][29] ),
    .S1(net1287),
    .X(_03371_));
 sg13g2_mux4_1 _09355_ (.S0(net1344),
    .A0(\dp.rf.rf[28][29] ),
    .A1(\dp.rf.rf[29][29] ),
    .A2(\dp.rf.rf[30][29] ),
    .A3(\dp.rf.rf[31][29] ),
    .S1(net1290),
    .X(_03372_));
 sg13g2_mux4_1 _09356_ (.S0(net1335),
    .A0(\dp.rf.rf[20][29] ),
    .A1(\dp.rf.rf[21][29] ),
    .A2(\dp.rf.rf[22][29] ),
    .A3(\dp.rf.rf[23][29] ),
    .S1(net1287),
    .X(_03373_));
 sg13g2_mux4_1 _09357_ (.S0(net1046),
    .A0(_03370_),
    .A1(_03371_),
    .A2(_03372_),
    .A3(_03373_),
    .S1(net1275),
    .X(_03374_));
 sg13g2_and2_1 _09358_ (.A(net1259),
    .B(_03374_),
    .X(_03375_));
 sg13g2_a22oi_1 _09359_ (.Y(_03376_),
    .B1(_03369_),
    .B2(_03375_),
    .A2(_03364_),
    .A1(net1050));
 sg13g2_buf_2 fanout993 (.A(_03749_),
    .X(net993));
 sg13g2_nor2_1 _09361_ (.A(net913),
    .B(_03376_),
    .Y(net154));
 sg13g2_mux4_1 _09362_ (.S0(net1337),
    .A0(\dp.rf.rf[8][30] ),
    .A1(\dp.rf.rf[9][30] ),
    .A2(\dp.rf.rf[10][30] ),
    .A3(\dp.rf.rf[11][30] ),
    .S1(net1288),
    .X(_03378_));
 sg13g2_mux4_1 _09363_ (.S0(net1337),
    .A0(\dp.rf.rf[0][30] ),
    .A1(\dp.rf.rf[1][30] ),
    .A2(\dp.rf.rf[2][30] ),
    .A3(\dp.rf.rf[3][30] ),
    .S1(net1288),
    .X(_03379_));
 sg13g2_mux4_1 _09364_ (.S0(net1338),
    .A0(\dp.rf.rf[12][30] ),
    .A1(\dp.rf.rf[13][30] ),
    .A2(\dp.rf.rf[14][30] ),
    .A3(\dp.rf.rf[15][30] ),
    .S1(net1289),
    .X(_03380_));
 sg13g2_mux4_1 _09365_ (.S0(net1338),
    .A0(\dp.rf.rf[4][30] ),
    .A1(\dp.rf.rf[5][30] ),
    .A2(\dp.rf.rf[6][30] ),
    .A3(\dp.rf.rf[7][30] ),
    .S1(net1289),
    .X(_03381_));
 sg13g2_mux4_1 _09366_ (.S0(net1046),
    .A0(_03378_),
    .A1(_03379_),
    .A2(_03380_),
    .A3(_03381_),
    .S1(net1276),
    .X(_03382_));
 sg13g2_mux4_1 _09367_ (.S0(net1338),
    .A0(\dp.rf.rf[24][30] ),
    .A1(\dp.rf.rf[25][30] ),
    .A2(\dp.rf.rf[26][30] ),
    .A3(\dp.rf.rf[27][30] ),
    .S1(net1289),
    .X(_03383_));
 sg13g2_mux4_1 _09368_ (.S0(net1338),
    .A0(\dp.rf.rf[16][30] ),
    .A1(\dp.rf.rf[17][30] ),
    .A2(\dp.rf.rf[18][30] ),
    .A3(\dp.rf.rf[19][30] ),
    .S1(net1289),
    .X(_03384_));
 sg13g2_mux4_1 _09369_ (.S0(net1338),
    .A0(\dp.rf.rf[28][30] ),
    .A1(\dp.rf.rf[29][30] ),
    .A2(\dp.rf.rf[30][30] ),
    .A3(\dp.rf.rf[31][30] ),
    .S1(net1289),
    .X(_03385_));
 sg13g2_mux4_1 _09370_ (.S0(net1338),
    .A0(\dp.rf.rf[20][30] ),
    .A1(\dp.rf.rf[21][30] ),
    .A2(\dp.rf.rf[22][30] ),
    .A3(\dp.rf.rf[23][30] ),
    .S1(net1289),
    .X(_03386_));
 sg13g2_mux4_1 _09371_ (.S0(net1046),
    .A0(_03383_),
    .A1(_03384_),
    .A2(_03385_),
    .A3(_03386_),
    .S1(net1276),
    .X(_03387_));
 sg13g2_and2_1 _09372_ (.A(net1259),
    .B(_03387_),
    .X(_03388_));
 sg13g2_a21oi_2 _09373_ (.B1(_03388_),
    .Y(_03389_),
    .A2(_03382_),
    .A1(_03307_));
 sg13g2_nor2_1 _09374_ (.A(net913),
    .B(_03389_),
    .Y(net156));
 sg13g2_nor2b_1 _09375_ (.A(net1319),
    .B_N(\dp.rf.rf[12][31] ),
    .Y(_03390_));
 sg13g2_a22oi_1 _09376_ (.Y(_03391_),
    .B1(net1086),
    .B2(_03390_),
    .A2(\dp.rf.rf[13][31] ),
    .A1(net1319));
 sg13g2_nor2b_1 _09377_ (.A(net1319),
    .B_N(\dp.rf.rf[14][31] ),
    .Y(_03392_));
 sg13g2_a22oi_1 _09378_ (.Y(_03393_),
    .B1(net1095),
    .B2(_03392_),
    .A2(\dp.rf.rf[15][31] ),
    .A1(net1319));
 sg13g2_nor2b_1 _09379_ (.A(net1315),
    .B_N(\dp.rf.rf[4][31] ),
    .Y(_03394_));
 sg13g2_a22oi_1 _09380_ (.Y(_03395_),
    .B1(net1080),
    .B2(_03394_),
    .A2(\dp.rf.rf[5][31] ),
    .A1(net1315));
 sg13g2_mux2_1 _09381_ (.A0(\dp.rf.rf[6][31] ),
    .A1(\dp.rf.rf[7][31] ),
    .S(net1319),
    .X(_03396_));
 sg13g2_o21ai_1 _09382_ (.B1(net1061),
    .Y(_03397_),
    .A1(net1074),
    .A2(_03396_));
 sg13g2_nor4_1 _09383_ (.A(_03391_),
    .B(_03393_),
    .C(_03395_),
    .D(_03397_),
    .Y(_03398_));
 sg13g2_nor2b_1 _09384_ (.A(net1319),
    .B_N(\dp.rf.rf[26][31] ),
    .Y(_03399_));
 sg13g2_a22oi_1 _09385_ (.Y(_03400_),
    .B1(net1095),
    .B2(_03399_),
    .A2(\dp.rf.rf[27][31] ),
    .A1(net1319));
 sg13g2_nor2b_1 _09386_ (.A(net1315),
    .B_N(\dp.rf.rf[24][31] ),
    .Y(_03401_));
 sg13g2_a22oi_1 _09387_ (.Y(_03402_),
    .B1(net1086),
    .B2(_03401_),
    .A2(\dp.rf.rf[25][31] ),
    .A1(net1315));
 sg13g2_nor2b_1 _09388_ (.A(net1315),
    .B_N(\dp.rf.rf[16][31] ),
    .Y(_03403_));
 sg13g2_a22oi_1 _09389_ (.Y(_03404_),
    .B1(net1080),
    .B2(_03403_),
    .A2(\dp.rf.rf[17][31] ),
    .A1(net1315));
 sg13g2_mux2_1 _09390_ (.A0(\dp.rf.rf[18][31] ),
    .A1(\dp.rf.rf[19][31] ),
    .S(net1318),
    .X(_03405_));
 sg13g2_o21ai_1 _09391_ (.B1(net1069),
    .Y(_03406_),
    .A1(net1074),
    .A2(_03405_));
 sg13g2_nor4_1 _09392_ (.A(_03400_),
    .B(_03402_),
    .C(_03404_),
    .D(_03406_),
    .Y(_03407_));
 sg13g2_nor2b_1 _09393_ (.A(net1321),
    .B_N(\dp.rf.rf[2][31] ),
    .Y(_03408_));
 sg13g2_a22oi_1 _09394_ (.Y(_03409_),
    .B1(net1074),
    .B2(_03408_),
    .A2(\dp.rf.rf[3][31] ),
    .A1(net1321));
 sg13g2_a21oi_1 _09395_ (.A1(net1316),
    .A2(\dp.rf.rf[1][31] ),
    .Y(_03410_),
    .B1(net1080));
 sg13g2_mux4_1 _09396_ (.S0(net1316),
    .A0(\dp.rf.rf[8][31] ),
    .A1(\dp.rf.rf[9][31] ),
    .A2(\dp.rf.rf[10][31] ),
    .A3(\dp.rf.rf[11][31] ),
    .S1(net1282),
    .X(_03411_));
 sg13g2_nor2_1 _09397_ (.A(net1045),
    .B(_03411_),
    .Y(_03412_));
 sg13g2_nor4_1 _09398_ (.A(net1105),
    .B(_03409_),
    .C(_03410_),
    .D(_03412_),
    .Y(_03413_));
 sg13g2_mux4_1 _09399_ (.S0(net1318),
    .A0(\dp.rf.rf[20][31] ),
    .A1(\dp.rf.rf[21][31] ),
    .A2(\dp.rf.rf[22][31] ),
    .A3(\dp.rf.rf[23][31] ),
    .S1(net1282),
    .X(_03414_));
 sg13g2_mux4_1 _09400_ (.S0(net1319),
    .A0(\dp.rf.rf[28][31] ),
    .A1(\dp.rf.rf[29][31] ),
    .A2(\dp.rf.rf[30][31] ),
    .A3(\dp.rf.rf[31][31] ),
    .S1(net1283),
    .X(_03415_));
 sg13g2_nor2b_1 _09401_ (.A(net1042),
    .B_N(_03415_),
    .Y(_03416_));
 sg13g2_a21o_1 _09402_ (.A2(_03414_),
    .A1(net951),
    .B1(_03416_),
    .X(_03417_));
 sg13g2_nor4_2 _09403_ (.A(_03398_),
    .B(_03407_),
    .C(_03413_),
    .Y(_03418_),
    .D(_03417_));
 sg13g2_buf_2 fanout992 (.A(_03756_),
    .X(net992));
 sg13g2_nor2_1 _09405_ (.A(net913),
    .B(_03418_),
    .Y(net157));
 sg13g2_nor2b_1 _09406_ (.A(net1349),
    .B_N(\dp.rf.rf[8][0] ),
    .Y(_03420_));
 sg13g2_a22oi_1 _09407_ (.Y(_03421_),
    .B1(net1090),
    .B2(_03420_),
    .A2(\dp.rf.rf[9][0] ),
    .A1(net1349));
 sg13g2_a21oi_1 _09408_ (.A1(net1356),
    .A2(\dp.rf.rf[1][0] ),
    .Y(_03422_),
    .B1(net1082));
 sg13g2_mux4_1 _09409_ (.S0(net1356),
    .A0(\dp.rf.rf[2][0] ),
    .A1(\dp.rf.rf[3][0] ),
    .A2(\dp.rf.rf[10][0] ),
    .A3(\dp.rf.rf[11][0] ),
    .S1(net1269),
    .X(_03423_));
 sg13g2_nor2_1 _09410_ (.A(net1102),
    .B(_03423_),
    .Y(_03424_));
 sg13g2_nor4_1 _09411_ (.A(net1103),
    .B(_03421_),
    .C(_03422_),
    .D(_03424_),
    .Y(_03425_));
 sg13g2_mux2_1 _09412_ (.A0(\dp.rf.rf[30][0] ),
    .A1(\dp.rf.rf[31][0] ),
    .S(net1328),
    .X(_03426_));
 sg13g2_nand2_1 _09413_ (.Y(_03427_),
    .A(_02663_),
    .B(_03426_));
 sg13g2_mux2_1 _09414_ (.A0(\dp.rf.rf[28][0] ),
    .A1(\dp.rf.rf[29][0] ),
    .S(net1328),
    .X(_03428_));
 sg13g2_nand3_1 _09415_ (.B(net1055),
    .C(_03428_),
    .A(net1067),
    .Y(_03429_));
 sg13g2_mux2_1 _09416_ (.A0(\dp.rf.rf[22][0] ),
    .A1(\dp.rf.rf[23][0] ),
    .S(net1356),
    .X(_03430_));
 sg13g2_nand3_1 _09417_ (.B(net1055),
    .C(_03430_),
    .A(net1052),
    .Y(_03431_));
 sg13g2_mux2_1 _09418_ (.A0(\dp.rf.rf[20][0] ),
    .A1(\dp.rf.rf[21][0] ),
    .S(net1356),
    .X(_03432_));
 sg13g2_nand3_1 _09419_ (.B(net1055),
    .C(_03432_),
    .A(net1059),
    .Y(_03433_));
 sg13g2_nand4_1 _09420_ (.B(_03429_),
    .C(_03431_),
    .A(_03427_),
    .Y(_03434_),
    .D(_03433_));
 sg13g2_nor2b_1 _09421_ (.A(net1327),
    .B_N(\dp.rf.rf[18][0] ),
    .Y(_03435_));
 sg13g2_a22oi_1 _09422_ (.Y(_03436_),
    .B1(net1074),
    .B2(_03435_),
    .A2(\dp.rf.rf[19][0] ),
    .A1(net1327));
 sg13g2_nor2b_1 _09423_ (.A(net1356),
    .B_N(\dp.rf.rf[16][0] ),
    .Y(_03437_));
 sg13g2_a22oi_1 _09424_ (.Y(_03438_),
    .B1(net1082),
    .B2(_03437_),
    .A2(\dp.rf.rf[17][0] ),
    .A1(net1355));
 sg13g2_nor2b_1 _09425_ (.A(net1355),
    .B_N(\dp.rf.rf[26][0] ),
    .Y(_03439_));
 sg13g2_a22oi_1 _09426_ (.Y(_03440_),
    .B1(net1097),
    .B2(_03439_),
    .A2(\dp.rf.rf[27][0] ),
    .A1(net1355));
 sg13g2_mux2_1 _09427_ (.A0(\dp.rf.rf[24][0] ),
    .A1(\dp.rf.rf[25][0] ),
    .S(net1355),
    .X(_03441_));
 sg13g2_o21ai_1 _09428_ (.B1(net1069),
    .Y(_03442_),
    .A1(net1090),
    .A2(_03441_));
 sg13g2_nor4_1 _09429_ (.A(_03436_),
    .B(_03438_),
    .C(_03440_),
    .D(_03442_),
    .Y(_03443_));
 sg13g2_mux4_1 _09430_ (.S0(net1356),
    .A0(\dp.rf.rf[4][0] ),
    .A1(\dp.rf.rf[5][0] ),
    .A2(\dp.rf.rf[6][0] ),
    .A3(\dp.rf.rf[7][0] ),
    .S1(net1291),
    .X(_03444_));
 sg13g2_mux4_1 _09431_ (.S0(net1356),
    .A0(\dp.rf.rf[12][0] ),
    .A1(\dp.rf.rf[13][0] ),
    .A2(\dp.rf.rf[14][0] ),
    .A3(\dp.rf.rf[15][0] ),
    .S1(net1291),
    .X(_03445_));
 sg13g2_nor2b_1 _09432_ (.A(_02815_),
    .B_N(_03445_),
    .Y(_03446_));
 sg13g2_a21o_1 _09433_ (.A2(_03444_),
    .A1(_02748_),
    .B1(_03446_),
    .X(_03447_));
 sg13g2_nor4_2 _09434_ (.A(_03425_),
    .B(_03434_),
    .C(_03443_),
    .Y(_03448_),
    .D(_03447_));
 sg13g2_inv_1 _09435_ (.Y(net133),
    .A(_03448_));
 sg13g2_mux4_1 _09436_ (.S0(net1380),
    .A0(\dp.rf.rf[20][1] ),
    .A1(\dp.rf.rf[21][1] ),
    .A2(\dp.rf.rf[22][1] ),
    .A3(\dp.rf.rf[23][1] ),
    .S1(net1298),
    .X(_03449_));
 sg13g2_mux4_1 _09437_ (.S0(net1380),
    .A0(\dp.rf.rf[28][1] ),
    .A1(\dp.rf.rf[29][1] ),
    .A2(\dp.rf.rf[30][1] ),
    .A3(\dp.rf.rf[31][1] ),
    .S1(net1298),
    .X(_03450_));
 sg13g2_nor2b_1 _09438_ (.A(net1043),
    .B_N(_03450_),
    .Y(_03451_));
 sg13g2_a21oi_1 _09439_ (.A1(net952),
    .A2(_03449_),
    .Y(_03452_),
    .B1(_03451_));
 sg13g2_mux2_1 _09440_ (.A0(\dp.rf.rf[1][1] ),
    .A1(\dp.rf.rf[9][1] ),
    .S(net1271),
    .X(_03453_));
 sg13g2_a221oi_1 _09441_ (.B2(net1377),
    .C1(net1297),
    .B1(_03453_),
    .A1(\dp.rf.rf[8][1] ),
    .Y(_03454_),
    .A2(_02731_));
 sg13g2_nor2b_1 _09442_ (.A(net1271),
    .B_N(\dp.rf.rf[2][1] ),
    .Y(_03455_));
 sg13g2_a22oi_1 _09443_ (.Y(_03456_),
    .B1(_02801_),
    .B2(_03455_),
    .A2(\dp.rf.rf[10][1] ),
    .A1(net1271));
 sg13g2_nor2b_1 _09444_ (.A(net1271),
    .B_N(\dp.rf.rf[3][1] ),
    .Y(_03457_));
 sg13g2_a22oi_1 _09445_ (.Y(_03458_),
    .B1(_02805_),
    .B2(_03457_),
    .A2(\dp.rf.rf[11][1] ),
    .A1(net1271));
 sg13g2_or4_1 _09446_ (.A(net1104),
    .B(_03454_),
    .C(_03456_),
    .D(_03458_),
    .X(_03459_));
 sg13g2_mux4_1 _09447_ (.S0(net1379),
    .A0(\dp.rf.rf[12][1] ),
    .A1(\dp.rf.rf[13][1] ),
    .A2(\dp.rf.rf[14][1] ),
    .A3(\dp.rf.rf[15][1] ),
    .S1(net1298),
    .X(_03460_));
 sg13g2_mux4_1 _09448_ (.S0(net1379),
    .A0(\dp.rf.rf[4][1] ),
    .A1(\dp.rf.rf[5][1] ),
    .A2(\dp.rf.rf[6][1] ),
    .A3(\dp.rf.rf[7][1] ),
    .S1(net1298),
    .X(_03461_));
 sg13g2_mux2_1 _09449_ (.A0(_03460_),
    .A1(_03461_),
    .S(net1048),
    .X(_03462_));
 sg13g2_nand2_1 _09450_ (.Y(_03463_),
    .A(net1064),
    .B(_03462_));
 sg13g2_nor2b_1 _09451_ (.A(net1378),
    .B_N(\dp.rf.rf[18][1] ),
    .Y(_03464_));
 sg13g2_a22oi_1 _09452_ (.Y(_03465_),
    .B1(net1077),
    .B2(_03464_),
    .A2(\dp.rf.rf[19][1] ),
    .A1(net1378));
 sg13g2_nor2b_1 _09453_ (.A(net1381),
    .B_N(\dp.rf.rf[16][1] ),
    .Y(_03466_));
 sg13g2_a22oi_1 _09454_ (.Y(_03467_),
    .B1(net1084),
    .B2(_03466_),
    .A2(\dp.rf.rf[17][1] ),
    .A1(net1381));
 sg13g2_nor2b_1 _09455_ (.A(net1380),
    .B_N(\dp.rf.rf[26][1] ),
    .Y(_03468_));
 sg13g2_a22oi_1 _09456_ (.Y(_03469_),
    .B1(net1098),
    .B2(_03468_),
    .A2(\dp.rf.rf[27][1] ),
    .A1(net1380));
 sg13g2_mux2_1 _09457_ (.A0(\dp.rf.rf[24][1] ),
    .A1(\dp.rf.rf[25][1] ),
    .S(net1381),
    .X(_03470_));
 sg13g2_o21ai_1 _09458_ (.B1(net1071),
    .Y(_03471_),
    .A1(net1092),
    .A2(_03470_));
 sg13g2_or4_1 _09459_ (.A(_03465_),
    .B(_03467_),
    .C(_03469_),
    .D(_03471_),
    .X(_03472_));
 sg13g2_nand4_1 _09460_ (.B(_03459_),
    .C(_03463_),
    .A(_03452_),
    .Y(net144),
    .D(_03472_));
 sg13g2_buf_2 fanout991 (.A(net992),
    .X(net991));
 sg13g2_mux2_1 _09462_ (.A0(\dp.rf.rf[2][2] ),
    .A1(\dp.rf.rf[3][2] ),
    .S(net1388),
    .X(_03474_));
 sg13g2_a221oi_1 _09463_ (.B2(net1299),
    .C1(net1272),
    .B1(_03474_),
    .A1(\dp.rf.rf[1][2] ),
    .Y(_03475_),
    .A2(_03097_));
 sg13g2_mux4_1 _09464_ (.S0(net1377),
    .A0(\dp.rf.rf[8][2] ),
    .A1(\dp.rf.rf[9][2] ),
    .A2(\dp.rf.rf[10][2] ),
    .A3(\dp.rf.rf[11][2] ),
    .S1(net1297),
    .X(_03476_));
 sg13g2_o21ai_1 _09465_ (.B1(net1050),
    .Y(_03477_),
    .A1(net1048),
    .A2(_03476_));
 sg13g2_or2_1 _09466_ (.X(_03478_),
    .B(_03477_),
    .A(_03475_));
 sg13g2_nor2b_1 _09467_ (.A(net1386),
    .B_N(\dp.rf.rf[22][2] ),
    .Y(_03479_));
 sg13g2_a22oi_1 _09468_ (.Y(_03480_),
    .B1(net1077),
    .B2(_03479_),
    .A2(\dp.rf.rf[23][2] ),
    .A1(net1386));
 sg13g2_nor2b_1 _09469_ (.A(net1386),
    .B_N(\dp.rf.rf[20][2] ),
    .Y(_03481_));
 sg13g2_a22oi_1 _09470_ (.Y(_03482_),
    .B1(net1084),
    .B2(_03481_),
    .A2(\dp.rf.rf[21][2] ),
    .A1(net1383));
 sg13g2_nor2b_1 _09471_ (.A(net1382),
    .B_N(\dp.rf.rf[30][2] ),
    .Y(_03483_));
 sg13g2_a22oi_1 _09472_ (.Y(_03484_),
    .B1(net1098),
    .B2(_03483_),
    .A2(\dp.rf.rf[31][2] ),
    .A1(net1383));
 sg13g2_mux2_1 _09473_ (.A0(\dp.rf.rf[28][2] ),
    .A1(\dp.rf.rf[29][2] ),
    .S(net1380),
    .X(_03485_));
 sg13g2_o21ai_1 _09474_ (.B1(net1057),
    .Y(_03486_),
    .A1(net1093),
    .A2(_03485_));
 sg13g2_or4_1 _09475_ (.A(_03480_),
    .B(_03482_),
    .C(_03484_),
    .D(_03486_),
    .X(_03487_));
 sg13g2_nor2b_1 _09476_ (.A(net1384),
    .B_N(\dp.rf.rf[26][2] ),
    .Y(_03488_));
 sg13g2_a22oi_1 _09477_ (.Y(_03489_),
    .B1(net1098),
    .B2(_03488_),
    .A2(\dp.rf.rf[27][2] ),
    .A1(net1384));
 sg13g2_nor2b_1 _09478_ (.A(net1382),
    .B_N(\dp.rf.rf[24][2] ),
    .Y(_03490_));
 sg13g2_a22oi_1 _09479_ (.Y(_03491_),
    .B1(net1092),
    .B2(_03490_),
    .A2(\dp.rf.rf[25][2] ),
    .A1(net1382));
 sg13g2_nor2b_1 _09480_ (.A(net1385),
    .B_N(\dp.rf.rf[16][2] ),
    .Y(_03492_));
 sg13g2_a22oi_1 _09481_ (.Y(_03493_),
    .B1(net1084),
    .B2(_03492_),
    .A2(\dp.rf.rf[17][2] ),
    .A1(net1385));
 sg13g2_mux2_1 _09482_ (.A0(\dp.rf.rf[18][2] ),
    .A1(\dp.rf.rf[19][2] ),
    .S(net1385),
    .X(_03494_));
 sg13g2_o21ai_1 _09483_ (.B1(net1071),
    .Y(_03495_),
    .A1(net1077),
    .A2(_03494_));
 sg13g2_or4_1 _09484_ (.A(_03489_),
    .B(_03491_),
    .C(_03493_),
    .D(_03495_),
    .X(_03496_));
 sg13g2_mux4_1 _09485_ (.S0(net1380),
    .A0(\dp.rf.rf[4][2] ),
    .A1(\dp.rf.rf[5][2] ),
    .A2(\dp.rf.rf[6][2] ),
    .A3(\dp.rf.rf[7][2] ),
    .S1(net1298),
    .X(_03497_));
 sg13g2_mux4_1 _09486_ (.S0(net1380),
    .A0(\dp.rf.rf[12][2] ),
    .A1(\dp.rf.rf[13][2] ),
    .A2(\dp.rf.rf[14][2] ),
    .A3(\dp.rf.rf[15][2] ),
    .S1(net1298),
    .X(_03498_));
 sg13g2_nor2b_1 _09487_ (.A(_02815_),
    .B_N(_03498_),
    .Y(_03499_));
 sg13g2_a21oi_1 _09488_ (.A1(_02748_),
    .A2(_03497_),
    .Y(_03500_),
    .B1(_03499_));
 sg13g2_and4_1 _09489_ (.A(_03478_),
    .B(_03487_),
    .C(_03496_),
    .D(_03500_),
    .X(_03501_));
 sg13g2_buf_4 fanout990 (.X(net990),
    .A(_03767_));
 sg13g2_inv_2 _09491_ (.Y(net155),
    .A(_03501_));
 sg13g2_nor2b_1 _09492_ (.A(net1260),
    .B_N(net1299),
    .Y(_03503_));
 sg13g2_mux2_1 _09493_ (.A0(\dp.rf.rf[6][3] ),
    .A1(\dp.rf.rf[7][3] ),
    .S(net1386),
    .X(_03504_));
 sg13g2_nand3_1 _09494_ (.B(_03503_),
    .C(_03504_),
    .A(net1049),
    .Y(_03505_));
 sg13g2_nor2_1 _09495_ (.A(net1260),
    .B(net1299),
    .Y(_03506_));
 sg13g2_mux2_1 _09496_ (.A0(\dp.rf.rf[4][3] ),
    .A1(\dp.rf.rf[5][3] ),
    .S(net1383),
    .X(_03507_));
 sg13g2_nand3_1 _09497_ (.B(_03506_),
    .C(_03507_),
    .A(net1049),
    .Y(_03508_));
 sg13g2_mux2_1 _09498_ (.A0(\dp.rf.rf[30][3] ),
    .A1(\dp.rf.rf[31][3] ),
    .S(net1383),
    .X(_03509_));
 sg13g2_nand4_1 _09499_ (.B(net1299),
    .C(net1272),
    .A(net1260),
    .Y(_03510_),
    .D(_03509_));
 sg13g2_nor2b_1 _09500_ (.A(net1299),
    .B_N(net1261),
    .Y(_03511_));
 sg13g2_mux2_1 _09501_ (.A0(\dp.rf.rf[28][3] ),
    .A1(\dp.rf.rf[29][3] ),
    .S(net1383),
    .X(_03512_));
 sg13g2_nand3_1 _09502_ (.B(_03511_),
    .C(_03512_),
    .A(net1272),
    .Y(_03513_));
 sg13g2_and4_1 _09503_ (.A(_03505_),
    .B(_03508_),
    .C(_03510_),
    .D(_03513_),
    .X(_03514_));
 sg13g2_mux2_1 _09504_ (.A0(\dp.rf.rf[14][3] ),
    .A1(\dp.rf.rf[15][3] ),
    .S(net1386),
    .X(_03515_));
 sg13g2_nand3_1 _09505_ (.B(_03503_),
    .C(_03515_),
    .A(net1272),
    .Y(_03516_));
 sg13g2_mux2_1 _09506_ (.A0(\dp.rf.rf[12][3] ),
    .A1(\dp.rf.rf[13][3] ),
    .S(net1388),
    .X(_03517_));
 sg13g2_nand3_1 _09507_ (.B(_03506_),
    .C(_03517_),
    .A(net1272),
    .Y(_03518_));
 sg13g2_mux2_1 _09508_ (.A0(\dp.rf.rf[22][3] ),
    .A1(\dp.rf.rf[23][3] ),
    .S(net1386),
    .X(_03519_));
 sg13g2_nand4_1 _09509_ (.B(net1300),
    .C(net1048),
    .A(net1261),
    .Y(_03520_),
    .D(_03519_));
 sg13g2_mux2_1 _09510_ (.A0(\dp.rf.rf[20][3] ),
    .A1(\dp.rf.rf[21][3] ),
    .S(net1386),
    .X(_03521_));
 sg13g2_nand3_1 _09511_ (.B(_03511_),
    .C(_03521_),
    .A(net1048),
    .Y(_03522_));
 sg13g2_and4_1 _09512_ (.A(_03516_),
    .B(_03518_),
    .C(_03520_),
    .D(_03522_),
    .X(_03523_));
 sg13g2_a21oi_1 _09513_ (.A1(_03514_),
    .A2(_03523_),
    .Y(_03524_),
    .B1(_03127_));
 sg13g2_nor2b_1 _09514_ (.A(net1388),
    .B_N(\dp.rf.rf[8][3] ),
    .Y(_03525_));
 sg13g2_a22oi_1 _09515_ (.Y(_03526_),
    .B1(net1092),
    .B2(_03525_),
    .A2(\dp.rf.rf[9][3] ),
    .A1(net1388));
 sg13g2_nor2b_1 _09516_ (.A(net1388),
    .B_N(\dp.rf.rf[10][3] ),
    .Y(_03527_));
 sg13g2_a22oi_1 _09517_ (.Y(_03528_),
    .B1(net1098),
    .B2(_03527_),
    .A2(\dp.rf.rf[11][3] ),
    .A1(net1388));
 sg13g2_mux2_1 _09518_ (.A0(\dp.rf.rf[2][3] ),
    .A1(\dp.rf.rf[3][3] ),
    .S(net1388),
    .X(_03529_));
 sg13g2_a221oi_1 _09519_ (.B2(net1299),
    .C1(net1274),
    .B1(_03529_),
    .A1(\dp.rf.rf[1][3] ),
    .Y(_03530_),
    .A2(_03097_));
 sg13g2_nor4_1 _09520_ (.A(net1103),
    .B(_03526_),
    .C(_03528_),
    .D(_03530_),
    .Y(_03531_));
 sg13g2_nor2b_1 _09521_ (.A(net1384),
    .B_N(\dp.rf.rf[26][3] ),
    .Y(_03532_));
 sg13g2_a22oi_1 _09522_ (.Y(_03533_),
    .B1(net1098),
    .B2(_03532_),
    .A2(\dp.rf.rf[27][3] ),
    .A1(net1384));
 sg13g2_nor2b_1 _09523_ (.A(net1382),
    .B_N(\dp.rf.rf[24][3] ),
    .Y(_03534_));
 sg13g2_a22oi_1 _09524_ (.Y(_03535_),
    .B1(net1092),
    .B2(_03534_),
    .A2(\dp.rf.rf[25][3] ),
    .A1(net1383));
 sg13g2_nor2b_1 _09525_ (.A(net1385),
    .B_N(\dp.rf.rf[18][3] ),
    .Y(_03536_));
 sg13g2_a22oi_1 _09526_ (.Y(_03537_),
    .B1(net1078),
    .B2(_03536_),
    .A2(\dp.rf.rf[19][3] ),
    .A1(net1384));
 sg13g2_mux2_1 _09527_ (.A0(\dp.rf.rf[16][3] ),
    .A1(\dp.rf.rf[17][3] ),
    .S(net1384),
    .X(_03538_));
 sg13g2_o21ai_1 _09528_ (.B1(net1071),
    .Y(_03539_),
    .A1(net1084),
    .A2(_03538_));
 sg13g2_nor4_1 _09529_ (.A(_03533_),
    .B(_03535_),
    .C(_03537_),
    .D(_03539_),
    .Y(_03540_));
 sg13g2_or2_1 _09530_ (.X(_03541_),
    .B(_03540_),
    .A(_03531_));
 sg13g2_buf_1 fanout989 (.A(_03771_),
    .X(net989));
 sg13g2_nor2_2 _09532_ (.A(_03524_),
    .B(_03541_),
    .Y(_03543_));
 sg13g2_inv_1 _09533_ (.Y(net158),
    .A(_03543_));
 sg13g2_mux4_1 _09534_ (.S0(net1355),
    .A0(\dp.rf.rf[8][4] ),
    .A1(\dp.rf.rf[9][4] ),
    .A2(\dp.rf.rf[10][4] ),
    .A3(\dp.rf.rf[11][4] ),
    .S1(net1291),
    .X(_03544_));
 sg13g2_mux4_1 _09535_ (.S0(net1357),
    .A0(\dp.rf.rf[0][4] ),
    .A1(\dp.rf.rf[1][4] ),
    .A2(\dp.rf.rf[2][4] ),
    .A3(\dp.rf.rf[3][4] ),
    .S1(net1291),
    .X(_03545_));
 sg13g2_mux2_1 _09536_ (.A0(_03544_),
    .A1(_03545_),
    .S(net1048),
    .X(_03546_));
 sg13g2_nand2_1 _09537_ (.Y(_03547_),
    .A(_02593_),
    .B(_03546_));
 sg13g2_nand3b_1 _09538_ (.B(net1277),
    .C(net1260),
    .Y(_03548_),
    .A_N(net1273));
 sg13g2_mux4_1 _09539_ (.S0(net1342),
    .A0(\dp.rf.rf[20][4] ),
    .A1(\dp.rf.rf[21][4] ),
    .A2(\dp.rf.rf[22][4] ),
    .A3(\dp.rf.rf[23][4] ),
    .S1(net1290),
    .X(_03549_));
 sg13g2_nor2b_1 _09540_ (.A(_03548_),
    .B_N(_03549_),
    .Y(_03550_));
 sg13g2_nor2b_1 _09541_ (.A(net1327),
    .B_N(\dp.rf.rf[18][4] ),
    .Y(_03551_));
 sg13g2_a22oi_1 _09542_ (.Y(_03552_),
    .B1(net1075),
    .B2(_03551_),
    .A2(\dp.rf.rf[19][4] ),
    .A1(net1343));
 sg13g2_nor2b_1 _09543_ (.A(net1327),
    .B_N(\dp.rf.rf[16][4] ),
    .Y(_03553_));
 sg13g2_a22oi_1 _09544_ (.Y(_03554_),
    .B1(net1081),
    .B2(_03553_),
    .A2(\dp.rf.rf[17][4] ),
    .A1(net1343));
 sg13g2_nor2b_1 _09545_ (.A(net1343),
    .B_N(\dp.rf.rf[26][4] ),
    .Y(_03555_));
 sg13g2_a22oi_1 _09546_ (.Y(_03556_),
    .B1(net1100),
    .B2(_03555_),
    .A2(\dp.rf.rf[27][4] ),
    .A1(net1343));
 sg13g2_mux2_1 _09547_ (.A0(\dp.rf.rf[24][4] ),
    .A1(\dp.rf.rf[25][4] ),
    .S(net1327),
    .X(_03557_));
 sg13g2_o21ai_1 _09548_ (.B1(net1072),
    .Y(_03558_),
    .A1(net1088),
    .A2(_03557_));
 sg13g2_nor4_1 _09549_ (.A(_03552_),
    .B(_03554_),
    .C(_03556_),
    .D(_03558_),
    .Y(_03559_));
 sg13g2_nor2b_1 _09550_ (.A(net1342),
    .B_N(\dp.rf.rf[30][4] ),
    .Y(_03560_));
 sg13g2_a21oi_1 _09551_ (.A1(net1344),
    .A2(\dp.rf.rf[31][4] ),
    .Y(_03561_),
    .B1(_03560_));
 sg13g2_mux2_1 _09552_ (.A0(\dp.rf.rf[28][4] ),
    .A1(\dp.rf.rf[29][4] ),
    .S(net1343),
    .X(_03562_));
 sg13g2_nand3_1 _09553_ (.B(net1054),
    .C(_03562_),
    .A(net1067),
    .Y(_03563_));
 sg13g2_o21ai_1 _09554_ (.B1(_03563_),
    .Y(_03564_),
    .A1(_02822_),
    .A2(_03561_));
 sg13g2_mux2_1 _09555_ (.A0(\dp.rf.rf[12][4] ),
    .A1(\dp.rf.rf[13][4] ),
    .S(net1327),
    .X(_03565_));
 sg13g2_nand3_1 _09556_ (.B(net1063),
    .C(_03565_),
    .A(net1067),
    .Y(_03566_));
 sg13g2_mux2_1 _09557_ (.A0(\dp.rf.rf[14][4] ),
    .A1(\dp.rf.rf[15][4] ),
    .S(net1355),
    .X(_03567_));
 sg13g2_nand3_1 _09558_ (.B(net1063),
    .C(_03567_),
    .A(_02642_),
    .Y(_03568_));
 sg13g2_mux2_1 _09559_ (.A0(\dp.rf.rf[4][4] ),
    .A1(\dp.rf.rf[5][4] ),
    .S(net1328),
    .X(_03569_));
 sg13g2_nand3_1 _09560_ (.B(net1063),
    .C(_03569_),
    .A(net1060),
    .Y(_03570_));
 sg13g2_mux2_1 _09561_ (.A0(\dp.rf.rf[6][4] ),
    .A1(\dp.rf.rf[7][4] ),
    .S(net1328),
    .X(_03571_));
 sg13g2_nand3_1 _09562_ (.B(net1061),
    .C(_03571_),
    .A(net1053),
    .Y(_03572_));
 sg13g2_nand4_1 _09563_ (.B(_03568_),
    .C(_03570_),
    .A(_03566_),
    .Y(_03573_),
    .D(_03572_));
 sg13g2_nor4_2 _09564_ (.A(_03550_),
    .B(_03559_),
    .C(_03564_),
    .Y(_03574_),
    .D(_03573_));
 sg13g2_nand2_2 _09565_ (.Y(net159),
    .A(_03547_),
    .B(_03574_));
 sg13g2_mux4_1 _09566_ (.S0(net1364),
    .A0(\dp.rf.rf[2][5] ),
    .A1(\dp.rf.rf[3][5] ),
    .A2(\dp.rf.rf[10][5] ),
    .A3(\dp.rf.rf[11][5] ),
    .S1(net1268),
    .X(_03575_));
 sg13g2_mux4_1 _09567_ (.S0(net1364),
    .A0(\dp.rf.rf[0][5] ),
    .A1(\dp.rf.rf[1][5] ),
    .A2(\dp.rf.rf[8][5] ),
    .A3(\dp.rf.rf[9][5] ),
    .S1(net1268),
    .X(_03576_));
 sg13g2_mux2_1 _09568_ (.A0(_03575_),
    .A1(_03576_),
    .S(net1102),
    .X(_03577_));
 sg13g2_mux4_1 _09569_ (.S0(net1368),
    .A0(\dp.rf.rf[4][5] ),
    .A1(\dp.rf.rf[5][5] ),
    .A2(\dp.rf.rf[6][5] ),
    .A3(\dp.rf.rf[7][5] ),
    .S1(net1295),
    .X(_03578_));
 sg13g2_mux4_1 _09570_ (.S0(net1368),
    .A0(\dp.rf.rf[20][5] ),
    .A1(\dp.rf.rf[21][5] ),
    .A2(\dp.rf.rf[22][5] ),
    .A3(\dp.rf.rf[23][5] ),
    .S1(net1295),
    .X(_03579_));
 sg13g2_nor2b_1 _09571_ (.A(_03548_),
    .B_N(_03579_),
    .Y(_03580_));
 sg13g2_a221oi_1 _09572_ (.B2(_02748_),
    .C1(_03580_),
    .B1(_03578_),
    .A1(net1051),
    .Y(_03581_),
    .A2(_03577_));
 sg13g2_mux4_1 _09573_ (.S0(net1368),
    .A0(\dp.rf.rf[24][5] ),
    .A1(\dp.rf.rf[25][5] ),
    .A2(\dp.rf.rf[26][5] ),
    .A3(\dp.rf.rf[27][5] ),
    .S1(net1295),
    .X(_03582_));
 sg13g2_mux4_1 _09574_ (.S0(net1368),
    .A0(\dp.rf.rf[16][5] ),
    .A1(\dp.rf.rf[17][5] ),
    .A2(\dp.rf.rf[18][5] ),
    .A3(\dp.rf.rf[19][5] ),
    .S1(net1295),
    .X(_03583_));
 sg13g2_mux2_1 _09575_ (.A0(_03582_),
    .A1(_03583_),
    .S(net1048),
    .X(_03584_));
 sg13g2_mux4_1 _09576_ (.S0(net1362),
    .A0(\dp.rf.rf[12][5] ),
    .A1(\dp.rf.rf[13][5] ),
    .A2(\dp.rf.rf[14][5] ),
    .A3(\dp.rf.rf[15][5] ),
    .S1(net1296),
    .X(_03585_));
 sg13g2_nor2b_1 _09577_ (.A(_02815_),
    .B_N(_03585_),
    .Y(_03586_));
 sg13g2_mux4_1 _09578_ (.S0(net1362),
    .A0(\dp.rf.rf[28][5] ),
    .A1(\dp.rf.rf[29][5] ),
    .A2(\dp.rf.rf[30][5] ),
    .A3(\dp.rf.rf[31][5] ),
    .S1(net1296),
    .X(_03587_));
 sg13g2_nor2b_1 _09579_ (.A(net1043),
    .B_N(_03587_),
    .Y(_03588_));
 sg13g2_a22oi_1 _09580_ (.Y(_03589_),
    .B1(_03586_),
    .B2(_03588_),
    .A2(_03584_),
    .A1(net1070));
 sg13g2_a21oi_2 _09581_ (.B1(net950),
    .Y(net160),
    .A2(_03589_),
    .A1(_03581_));
 sg13g2_nor2b_1 _09582_ (.A(net1362),
    .B_N(\dp.rf.rf[18][6] ),
    .Y(_03590_));
 sg13g2_a22oi_1 _09583_ (.Y(_03591_),
    .B1(net1076),
    .B2(_03590_),
    .A2(\dp.rf.rf[19][6] ),
    .A1(net1362));
 sg13g2_nor2b_1 _09584_ (.A(net1362),
    .B_N(\dp.rf.rf[16][6] ),
    .Y(_03592_));
 sg13g2_a22oi_1 _09585_ (.Y(_03593_),
    .B1(net1083),
    .B2(_03592_),
    .A2(\dp.rf.rf[17][6] ),
    .A1(net1362));
 sg13g2_nor2b_1 _09586_ (.A(net1362),
    .B_N(\dp.rf.rf[26][6] ),
    .Y(_03594_));
 sg13g2_a22oi_1 _09587_ (.Y(_03595_),
    .B1(net1099),
    .B2(_03594_),
    .A2(\dp.rf.rf[27][6] ),
    .A1(net1362));
 sg13g2_mux2_1 _09588_ (.A0(\dp.rf.rf[24][6] ),
    .A1(\dp.rf.rf[25][6] ),
    .S(net1363),
    .X(_03596_));
 sg13g2_o21ai_1 _09589_ (.B1(net1070),
    .Y(_03597_),
    .A1(net1091),
    .A2(_03596_));
 sg13g2_nor4_1 _09590_ (.A(_03591_),
    .B(_03593_),
    .C(_03595_),
    .D(_03597_),
    .Y(_03598_));
 sg13g2_mux4_1 _09591_ (.S0(net1363),
    .A0(\dp.rf.rf[20][6] ),
    .A1(\dp.rf.rf[21][6] ),
    .A2(\dp.rf.rf[22][6] ),
    .A3(\dp.rf.rf[23][6] ),
    .S1(net1294),
    .X(_03599_));
 sg13g2_mux4_1 _09592_ (.S0(net1363),
    .A0(\dp.rf.rf[28][6] ),
    .A1(\dp.rf.rf[29][6] ),
    .A2(\dp.rf.rf[30][6] ),
    .A3(\dp.rf.rf[31][6] ),
    .S1(net1294),
    .X(_03600_));
 sg13g2_nor2b_1 _09593_ (.A(net1043),
    .B_N(_03600_),
    .Y(_03601_));
 sg13g2_a21o_1 _09594_ (.A2(_03599_),
    .A1(net952),
    .B1(_03601_),
    .X(_03602_));
 sg13g2_mux4_1 _09595_ (.S0(net1361),
    .A0(\dp.rf.rf[2][6] ),
    .A1(\dp.rf.rf[3][6] ),
    .A2(\dp.rf.rf[10][6] ),
    .A3(\dp.rf.rf[11][6] ),
    .S1(net1267),
    .X(_03603_));
 sg13g2_inv_1 _09596_ (.Y(_03604_),
    .A(_03603_));
 sg13g2_mux2_1 _09597_ (.A0(\dp.rf.rf[1][6] ),
    .A1(\dp.rf.rf[9][6] ),
    .S(net1267),
    .X(_03605_));
 sg13g2_a221oi_1 _09598_ (.B2(net1361),
    .C1(net1293),
    .B1(_03605_),
    .A1(\dp.rf.rf[8][6] ),
    .Y(_03606_),
    .A2(_02731_));
 sg13g2_a22oi_1 _09599_ (.Y(_03607_),
    .B1(_03606_),
    .B2(net1103),
    .A2(_03604_),
    .A1(net1293));
 sg13g2_mux4_1 _09600_ (.S0(net1360),
    .A0(\dp.rf.rf[12][6] ),
    .A1(\dp.rf.rf[13][6] ),
    .A2(\dp.rf.rf[14][6] ),
    .A3(\dp.rf.rf[15][6] ),
    .S1(net1294),
    .X(_03608_));
 sg13g2_nand2_1 _09601_ (.Y(_03609_),
    .A(net1267),
    .B(_03608_));
 sg13g2_mux4_1 _09602_ (.S0(net1360),
    .A0(\dp.rf.rf[4][6] ),
    .A1(\dp.rf.rf[5][6] ),
    .A2(\dp.rf.rf[6][6] ),
    .A3(\dp.rf.rf[7][6] ),
    .S1(net1293),
    .X(_03610_));
 sg13g2_nand2_1 _09603_ (.Y(_03611_),
    .A(net1048),
    .B(_03610_));
 sg13g2_a21oi_1 _09604_ (.A1(_03609_),
    .A2(_03611_),
    .Y(_03612_),
    .B1(_02746_));
 sg13g2_nor4_2 _09605_ (.A(_03598_),
    .B(_03602_),
    .C(_03607_),
    .Y(_03613_),
    .D(_03612_));
 sg13g2_buf_2 fanout988 (.A(net989),
    .X(net988));
 sg13g2_inv_1 _09607_ (.Y(net161),
    .A(_03613_));
 sg13g2_nand2_1 _09608_ (.Y(_03615_),
    .A(net1357),
    .B(\dp.rf.rf[13][7] ));
 sg13g2_nand2b_1 _09609_ (.Y(_03616_),
    .B(\dp.rf.rf[12][7] ),
    .A_N(net1359));
 sg13g2_a21oi_1 _09610_ (.A1(_03615_),
    .A2(_03616_),
    .Y(_03617_),
    .B1(net1090));
 sg13g2_nand2_1 _09611_ (.Y(_03618_),
    .A(net1359),
    .B(\dp.rf.rf[15][7] ));
 sg13g2_nand2b_1 _09612_ (.Y(_03619_),
    .B(\dp.rf.rf[14][7] ),
    .A_N(net1359));
 sg13g2_a21oi_1 _09613_ (.A1(_03618_),
    .A2(_03619_),
    .Y(_03620_),
    .B1(net1097));
 sg13g2_o21ai_1 _09614_ (.B1(net1064),
    .Y(_03621_),
    .A1(_03617_),
    .A2(_03620_));
 sg13g2_mux4_1 _09615_ (.S0(net1358),
    .A0(\dp.rf.rf[8][7] ),
    .A1(\dp.rf.rf[9][7] ),
    .A2(\dp.rf.rf[10][7] ),
    .A3(\dp.rf.rf[11][7] ),
    .S1(net1291),
    .X(_03622_));
 sg13g2_nand2_1 _09616_ (.Y(_03623_),
    .A(net1269),
    .B(_03622_));
 sg13g2_mux4_1 _09617_ (.S0(net1358),
    .A0(\dp.rf.rf[0][7] ),
    .A1(\dp.rf.rf[1][7] ),
    .A2(\dp.rf.rf[2][7] ),
    .A3(\dp.rf.rf[3][7] ),
    .S1(net1292),
    .X(_03624_));
 sg13g2_nand2_1 _09618_ (.Y(_03625_),
    .A(net1048),
    .B(_03624_));
 sg13g2_a21oi_1 _09619_ (.A1(_03623_),
    .A2(_03625_),
    .Y(_03626_),
    .B1(_03215_));
 sg13g2_nor2b_1 _09620_ (.A(net1364),
    .B_N(\dp.rf.rf[26][7] ),
    .Y(_03627_));
 sg13g2_a22oi_1 _09621_ (.Y(_03628_),
    .B1(net1097),
    .B2(_03627_),
    .A2(\dp.rf.rf[27][7] ),
    .A1(net1364));
 sg13g2_nor2b_1 _09622_ (.A(net1365),
    .B_N(\dp.rf.rf[18][7] ),
    .Y(_03629_));
 sg13g2_a22oi_1 _09623_ (.Y(_03630_),
    .B1(net1078),
    .B2(_03629_),
    .A2(\dp.rf.rf[19][7] ),
    .A1(net1365));
 sg13g2_nor2b_1 _09624_ (.A(net1365),
    .B_N(\dp.rf.rf[24][7] ),
    .Y(_03631_));
 sg13g2_a22oi_1 _09625_ (.Y(_03632_),
    .B1(net1091),
    .B2(_03631_),
    .A2(\dp.rf.rf[25][7] ),
    .A1(net1365));
 sg13g2_mux2_1 _09626_ (.A0(\dp.rf.rf[16][7] ),
    .A1(\dp.rf.rf[17][7] ),
    .S(net1365),
    .X(_03633_));
 sg13g2_o21ai_1 _09627_ (.B1(net1070),
    .Y(_03634_),
    .A1(net1083),
    .A2(_03633_));
 sg13g2_nor4_1 _09628_ (.A(_03628_),
    .B(_03630_),
    .C(_03632_),
    .D(_03634_),
    .Y(_03635_));
 sg13g2_mux2_1 _09629_ (.A0(\dp.rf.rf[6][7] ),
    .A1(\dp.rf.rf[7][7] ),
    .S(net1358),
    .X(_03636_));
 sg13g2_nand3_1 _09630_ (.B(net1065),
    .C(_03636_),
    .A(net1052),
    .Y(_03637_));
 sg13g2_mux2_1 _09631_ (.A0(\dp.rf.rf[30][7] ),
    .A1(\dp.rf.rf[31][7] ),
    .S(net1364),
    .X(_03638_));
 sg13g2_nand2_1 _09632_ (.Y(_03639_),
    .A(_02663_),
    .B(_03638_));
 sg13g2_mux2_1 _09633_ (.A0(\dp.rf.rf[4][7] ),
    .A1(\dp.rf.rf[5][7] ),
    .S(net1358),
    .X(_03640_));
 sg13g2_nand3_1 _09634_ (.B(net1065),
    .C(_03640_),
    .A(net1059),
    .Y(_03641_));
 sg13g2_mux2_1 _09635_ (.A0(\dp.rf.rf[20][7] ),
    .A1(\dp.rf.rf[21][7] ),
    .S(net1364),
    .X(_03642_));
 sg13g2_nand3_1 _09636_ (.B(net1056),
    .C(_03642_),
    .A(net1059),
    .Y(_03643_));
 sg13g2_nand4_1 _09637_ (.B(_03639_),
    .C(_03641_),
    .A(_03637_),
    .Y(_03644_),
    .D(_03643_));
 sg13g2_mux2_1 _09638_ (.A0(\dp.rf.rf[28][7] ),
    .A1(\dp.rf.rf[29][7] ),
    .S(net1364),
    .X(_03645_));
 sg13g2_nand3_1 _09639_ (.B(net1057),
    .C(_03645_),
    .A(net1068),
    .Y(_03646_));
 sg13g2_mux2_1 _09640_ (.A0(\dp.rf.rf[22][7] ),
    .A1(\dp.rf.rf[23][7] ),
    .S(net1358),
    .X(_03647_));
 sg13g2_nand3_1 _09641_ (.B(net1056),
    .C(_03647_),
    .A(net1052),
    .Y(_03648_));
 sg13g2_nand2_1 _09642_ (.Y(_03649_),
    .A(_03646_),
    .B(_03648_));
 sg13g2_nor4_2 _09643_ (.A(_03626_),
    .B(_03635_),
    .C(_03644_),
    .Y(_03650_),
    .D(_03649_));
 sg13g2_nand2_2 _09644_ (.Y(net162),
    .A(_03621_),
    .B(_03650_));
 sg13g2_buf_4 fanout987 (.X(net987),
    .A(_03775_));
 sg13g2_buf_2 fanout986 (.A(_03799_),
    .X(net986));
 sg13g2_buf_2 fanout985 (.A(_03812_),
    .X(net985));
 sg13g2_nor2_1 _09648_ (.A(net1228),
    .B(net1114),
    .Y(_03654_));
 sg13g2_buf_1 fanout984 (.A(_03859_),
    .X(net984));
 sg13g2_buf_2 fanout983 (.A(_03859_),
    .X(net983));
 sg13g2_buf_2 fanout982 (.A(net983),
    .X(net982));
 sg13g2_buf_2 fanout981 (.A(_03917_),
    .X(net981));
 sg13g2_buf_2 fanout980 (.A(net981),
    .X(net980));
 sg13g2_buf_2 fanout979 (.A(net980),
    .X(net979));
 sg13g2_buf_2 fanout978 (.A(net980),
    .X(net978));
 sg13g2_nand3b_1 _09656_ (.B(net12),
    .C(net1),
    .Y(_03662_),
    .A_N(net1248));
 sg13g2_buf_4 fanout977 (.X(net977),
    .A(net981));
 sg13g2_buf_2 fanout976 (.A(net977),
    .X(net976));
 sg13g2_buf_1 fanout975 (.A(_03917_),
    .X(net975));
 sg13g2_nand3b_1 _09660_ (.B(net1255),
    .C(net27),
    .Y(_03666_),
    .A_N(net1252));
 sg13g2_buf_2 fanout974 (.A(net975),
    .X(net974));
 sg13g2_buf_2 fanout973 (.A(_03917_),
    .X(net973));
 sg13g2_buf_2 fanout972 (.A(net973),
    .X(net972));
 sg13g2_buf_2 fanout971 (.A(net973),
    .X(net971));
 sg13g2_buf_4 fanout970 (.X(net970),
    .A(net973));
 sg13g2_nor2b_1 _09666_ (.A(_00010_),
    .B_N(net1170),
    .Y(_03672_));
 sg13g2_o21ai_1 _09667_ (.B1(_03672_),
    .Y(_03673_),
    .A1(net1035),
    .A2(net1021));
 sg13g2_o21ai_1 _09668_ (.B1(_03673_),
    .Y(_03674_),
    .A1(net1170),
    .A2(_00008_));
 sg13g2_buf_2 fanout969 (.A(_03964_),
    .X(net969));
 sg13g2_nand2b_1 _09670_ (.Y(_03676_),
    .B(net1114),
    .A_N(net1228));
 sg13g2_buf_4 fanout968 (.X(net968),
    .A(_03973_));
 sg13g2_buf_2 fanout967 (.A(net968),
    .X(net967));
 sg13g2_buf_2 fanout966 (.A(net967),
    .X(net966));
 sg13g2_nor2b_1 _09674_ (.A(net1170),
    .B_N(_00012_),
    .Y(_03680_));
 sg13g2_a22oi_1 _09675_ (.Y(_03681_),
    .B1(net1007),
    .B2(_03680_),
    .A2(_00014_),
    .A1(net1170));
 sg13g2_buf_2 fanout965 (.A(_03980_),
    .X(net965));
 sg13g2_nand2_1 _09677_ (.Y(_03683_),
    .A(net1228),
    .B(net1114));
 sg13g2_buf_2 fanout964 (.A(net965),
    .X(net964));
 sg13g2_nor2b_1 _09679_ (.A(net1170),
    .B_N(_00013_),
    .Y(_03685_));
 sg13g2_a22oi_1 _09680_ (.Y(_03686_),
    .B1(net1006),
    .B2(_03685_),
    .A2(_00015_),
    .A1(net1170));
 sg13g2_buf_2 fanout963 (.A(net965),
    .X(net963));
 sg13g2_buf_2 fanout962 (.A(_04250_),
    .X(net962));
 sg13g2_nand2b_1 _09683_ (.Y(_03689_),
    .B(net1228),
    .A_N(net1114));
 sg13g2_buf_4 fanout961 (.X(net961),
    .A(_04250_));
 sg13g2_nor2b_1 _09685_ (.A(net1171),
    .B_N(_00009_),
    .Y(_03691_));
 sg13g2_a22oi_1 _09686_ (.Y(_03692_),
    .B1(net1004),
    .B2(_03691_),
    .A2(_00011_),
    .A1(net1171));
 sg13g2_or3_1 _09687_ (.A(_03681_),
    .B(_03686_),
    .C(_03692_),
    .X(_03693_));
 sg13g2_buf_2 fanout960 (.A(_04305_),
    .X(net960));
 sg13g2_buf_2 fanout959 (.A(net960),
    .X(net959));
 sg13g2_buf_2 fanout958 (.A(_04305_),
    .X(net958));
 sg13g2_nor2b_1 _09691_ (.A(net1393),
    .B_N(net1399),
    .Y(_03697_));
 sg13g2_o21ai_1 _09692_ (.B1(_03697_),
    .Y(_03698_),
    .A1(net1034),
    .A2(net1020));
 sg13g2_buf_2 fanout957 (.A(_01053_),
    .X(net957));
 sg13g2_buf_2 fanout956 (.A(net957),
    .X(net956));
 sg13g2_a22oi_1 _09695_ (.Y(_03701_),
    .B1(_03693_),
    .B2(net947),
    .A2(_03674_),
    .A1(net1040));
 sg13g2_o21ai_1 _09696_ (.B1(net1392),
    .Y(_03702_),
    .A1(net1025),
    .A2(net1011));
 sg13g2_buf_4 fanout955 (.X(net955),
    .A(net956));
 sg13g2_buf_4 fanout954 (.X(net954),
    .A(_01053_));
 sg13g2_nand2_1 _09699_ (.Y(_03705_),
    .A(net1144),
    .B(_00031_));
 sg13g2_buf_4 fanout953 (.X(net953),
    .A(net954));
 sg13g2_nand2b_1 _09701_ (.Y(_03707_),
    .B(_00029_),
    .A_N(net1144));
 sg13g2_buf_2 fanout952 (.A(_02770_),
    .X(net952));
 sg13g2_buf_2 fanout951 (.A(_02770_),
    .X(net951));
 sg13g2_buf_1 fanout950 (.A(_03304_),
    .X(net950));
 sg13g2_nand3_1 _09705_ (.B(net1110),
    .C(net1398),
    .A(net1217),
    .Y(_03711_));
 sg13g2_a21oi_1 _09706_ (.A1(_03705_),
    .A2(_03707_),
    .Y(_03712_),
    .B1(_03711_));
 sg13g2_nand2_1 _09707_ (.Y(_03713_),
    .A(net1144),
    .B(_00030_));
 sg13g2_nand2b_1 _09708_ (.Y(_03714_),
    .B(_00028_),
    .A_N(net1145));
 sg13g2_inv_1 _09709_ (.Y(_03715_),
    .A(net1396));
 sg13g2_a22oi_1 _09710_ (.Y(_03716_),
    .B1(net1003),
    .B2(net1008),
    .A2(_03714_),
    .A1(_03713_));
 sg13g2_nand2_1 _09711_ (.Y(_03717_),
    .A(net1146),
    .B(_00019_));
 sg13g2_buf_2 fanout949 (.A(net950),
    .X(net949));
 sg13g2_nand2b_1 _09713_ (.Y(_03719_),
    .B(_00017_),
    .A_N(net1172));
 sg13g2_buf_1 fanout948 (.A(_03698_),
    .X(net948));
 sg13g2_a22oi_1 _09715_ (.Y(_03721_),
    .B1(net1399),
    .B2(net1005),
    .A2(_03719_),
    .A1(_03717_));
 sg13g2_buf_2 fanout947 (.A(_03698_),
    .X(net947));
 sg13g2_nand2_1 _09717_ (.Y(_03723_),
    .A(net1172),
    .B(_00018_));
 sg13g2_nand2b_1 _09718_ (.Y(_03724_),
    .B(_00016_),
    .A_N(net1170));
 sg13g2_or2_2 _09719_ (.X(_03725_),
    .B(net1114),
    .A(net1227));
 sg13g2_buf_2 fanout946 (.A(_03702_),
    .X(net946));
 sg13g2_a22oi_1 _09721_ (.Y(_03727_),
    .B1(net1399),
    .B2(net998),
    .A2(_03724_),
    .A1(_03723_));
 sg13g2_nor4_1 _09722_ (.A(_03712_),
    .B(_03716_),
    .C(_03721_),
    .D(_03727_),
    .Y(_03728_));
 sg13g2_nor2_1 _09723_ (.A(net945),
    .B(_03728_),
    .Y(_03729_));
 sg13g2_or2_1 _09724_ (.X(_03730_),
    .B(net1016),
    .A(net1030));
 sg13g2_buf_2 fanout945 (.A(_03702_),
    .X(net945));
 sg13g2_buf_1 fanout944 (.A(_03730_),
    .X(net944));
 sg13g2_buf_2 fanout943 (.A(net944),
    .X(net943));
 sg13g2_inv_2 _09728_ (.Y(_03734_),
    .A(net1391));
 sg13g2_nand2b_2 _09729_ (.Y(_03735_),
    .B(net1106),
    .A_N(net1396));
 sg13g2_buf_2 fanout942 (.A(net944),
    .X(net942));
 sg13g2_nor2_2 _09731_ (.A(net995),
    .B(_03735_),
    .Y(_03737_));
 sg13g2_buf_1 fanout941 (.A(net944),
    .X(net941));
 sg13g2_buf_2 fanout940 (.A(net941),
    .X(net940));
 sg13g2_buf_2 fanout939 (.A(net941),
    .X(net939));
 sg13g2_mux4_1 _09735_ (.S0(net1170),
    .A0(_00020_),
    .A1(_00022_),
    .A2(_00021_),
    .A3(_00023_),
    .S1(net1226),
    .X(_03741_));
 sg13g2_nand3_1 _09736_ (.B(net925),
    .C(_03741_),
    .A(net936),
    .Y(_03742_));
 sg13g2_nor2_2 _09737_ (.A(net1216),
    .B(net1150),
    .Y(_03743_));
 sg13g2_buf_2 fanout938 (.A(net944),
    .X(net938));
 sg13g2_nor3_2 _09739_ (.A(net1113),
    .B(net1399),
    .C(net1393),
    .Y(_03745_));
 sg13g2_nand2_2 _09740_ (.Y(_03746_),
    .A(_03743_),
    .B(_03745_));
 sg13g2_and2_1 _09741_ (.A(net939),
    .B(_03746_),
    .X(_03747_));
 sg13g2_buf_2 fanout937 (.A(net938),
    .X(net937));
 sg13g2_and2_1 _09743_ (.A(net1399),
    .B(net1393),
    .X(_03749_));
 sg13g2_buf_1 fanout936 (.A(net938),
    .X(net936));
 sg13g2_mux2_1 _09745_ (.A0(_00024_),
    .A1(_00026_),
    .S(net1172),
    .X(_03751_));
 sg13g2_nand3_1 _09746_ (.B(_03749_),
    .C(_03751_),
    .A(net1040),
    .Y(_03752_));
 sg13g2_buf_2 fanout935 (.A(net938),
    .X(net935));
 sg13g2_buf_1 fanout934 (.A(_03730_),
    .X(net934));
 sg13g2_buf_2 fanout933 (.A(net934),
    .X(net933));
 sg13g2_nor2b_2 _09750_ (.A(net1106),
    .B_N(net1396),
    .Y(_03756_));
 sg13g2_buf_2 fanout932 (.A(net933),
    .X(net932));
 sg13g2_buf_2 fanout931 (.A(net932),
    .X(net931));
 sg13g2_mux2_1 _09753_ (.A0(_00025_),
    .A1(_00027_),
    .S(net1172),
    .X(_03759_));
 sg13g2_nand4_1 _09754_ (.B(net1393),
    .C(_03756_),
    .A(net1226),
    .Y(_03760_),
    .D(_03759_));
 sg13g2_nand4_1 _09755_ (.B(net912),
    .C(_03752_),
    .A(_03742_),
    .Y(_03761_),
    .D(_03760_));
 sg13g2_buf_1 fanout930 (.A(net934),
    .X(net930));
 sg13g2_buf_1 fanout929 (.A(net930),
    .X(net929));
 sg13g2_nor2b_1 _09758_ (.A(net1171),
    .B_N(_00004_),
    .Y(_03764_));
 sg13g2_a22oi_1 _09759_ (.Y(_03765_),
    .B1(net1007),
    .B2(_03764_),
    .A2(_00006_),
    .A1(net1171));
 sg13g2_buf_2 fanout928 (.A(net930),
    .X(net928));
 sg13g2_nand2b_1 _09761_ (.Y(_03767_),
    .B(net1229),
    .A_N(net1182));
 sg13g2_buf_1 fanout927 (.A(net930),
    .X(net927));
 sg13g2_nor2b_1 _09763_ (.A(net1112),
    .B_N(_00001_),
    .Y(_03769_));
 sg13g2_a22oi_1 _09764_ (.Y(_03770_),
    .B1(net990),
    .B2(_03769_),
    .A2(_00005_),
    .A1(net1112));
 sg13g2_or2_1 _09765_ (.X(_03771_),
    .B(net1394),
    .A(net1401));
 sg13g2_buf_2 fanout926 (.A(net930),
    .X(net926));
 sg13g2_buf_2 fanout925 (.A(_03737_),
    .X(net925));
 sg13g2_buf_2 fanout924 (.A(_03786_),
    .X(net924));
 sg13g2_nand2_2 _09769_ (.Y(_03775_),
    .A(net1229),
    .B(net1182));
 sg13g2_buf_2 fanout923 (.A(net924),
    .X(net923));
 sg13g2_buf_2 fanout922 (.A(net923),
    .X(net922));
 sg13g2_nor2b_1 _09772_ (.A(net1112),
    .B_N(_00003_),
    .Y(_03778_));
 sg13g2_a22oi_1 _09773_ (.Y(_03779_),
    .B1(_03775_),
    .B2(_03778_),
    .A2(_00007_),
    .A1(net1112));
 sg13g2_or4_1 _09774_ (.A(_03765_),
    .B(_03770_),
    .C(net989),
    .D(_03779_),
    .X(_03780_));
 sg13g2_or3_1 _09775_ (.A(net1214),
    .B(net1144),
    .C(net1108),
    .X(_03781_));
 sg13g2_buf_2 fanout921 (.A(net924),
    .X(net921));
 sg13g2_o21ai_1 _09777_ (.B1(_03781_),
    .Y(_03783_),
    .A1(net1035),
    .A2(net1021));
 sg13g2_buf_2 fanout920 (.A(net924),
    .X(net920));
 sg13g2_nor2b_1 _09779_ (.A(_00000_),
    .B_N(_03783_),
    .Y(_03785_));
 sg13g2_nor2_1 _09780_ (.A(net1037),
    .B(net1022),
    .Y(_03786_));
 sg13g2_buf_2 fanout919 (.A(net924),
    .X(net919));
 sg13g2_buf_2 fanout918 (.A(net924),
    .X(net918));
 sg13g2_buf_2 fanout917 (.A(_04457_),
    .X(net917));
 sg13g2_nand2_2 _09784_ (.Y(_03790_),
    .A(net1191),
    .B(net1041));
 sg13g2_buf_4 fanout916 (.X(net916),
    .A(_04457_));
 sg13g2_nor3_1 _09786_ (.A(_00002_),
    .B(net921),
    .C(_03790_),
    .Y(_03792_));
 sg13g2_a22oi_1 _09787_ (.Y(_03793_),
    .B1(_03785_),
    .B2(_03792_),
    .A2(_03780_),
    .A1(net935));
 sg13g2_nor4_1 _09788_ (.A(_03701_),
    .B(_03729_),
    .C(_03761_),
    .D(_03793_),
    .Y(_03794_));
 sg13g2_buf_2 fanout915 (.A(_04481_),
    .X(net915));
 sg13g2_inv_1 _09790_ (.Y(_03796_),
    .A(net27));
 sg13g2_buf_2 fanout914 (.A(net915),
    .X(net914));
 sg13g2_nor2_1 _09792_ (.A(_03796_),
    .B(net1249),
    .Y(_03798_));
 sg13g2_or2_1 _09793_ (.X(_03799_),
    .B(net1254),
    .A(net1251));
 sg13g2_buf_2 fanout913 (.A(_02976_),
    .X(net913));
 sg13g2_or2_1 _09795_ (.X(_03801_),
    .B(net1036),
    .A(_03799_));
 sg13g2_buf_2 fanout912 (.A(_03747_),
    .X(net912));
 sg13g2_buf_2 fanout911 (.A(_03831_),
    .X(net911));
 sg13g2_nor2b_1 _09798_ (.A(net1237),
    .B_N(net1241),
    .Y(_03804_));
 sg13g2_o21ai_1 _09799_ (.B1(_03804_),
    .Y(_03805_),
    .A1(_03798_),
    .A2(_03801_));
 sg13g2_nand2_1 _09800_ (.Y(_03806_),
    .A(net27),
    .B(net1249));
 sg13g2_buf_2 fanout910 (.A(_03831_),
    .X(net910));
 sg13g2_nor2b_1 _09802_ (.A(net1253),
    .B_N(net1239),
    .Y(_03808_));
 sg13g2_a21oi_1 _09803_ (.A1(net24),
    .A2(_02576_),
    .Y(_03809_),
    .B1(_03808_));
 sg13g2_or4_1 _09804_ (.A(net1237),
    .B(_03801_),
    .C(_03806_),
    .D(_03809_),
    .X(_03810_));
 sg13g2_buf_2 fanout909 (.A(net910),
    .X(net909));
 sg13g2_nand2b_1 _09806_ (.Y(_03812_),
    .B(net1249),
    .A_N(net27));
 sg13g2_buf_2 fanout908 (.A(net909),
    .X(net908));
 sg13g2_nand3_1 _09808_ (.B(net12),
    .C(net1248),
    .A(net1),
    .Y(_03814_));
 sg13g2_buf_2 fanout907 (.A(_03831_),
    .X(net907));
 sg13g2_nor3_1 _09810_ (.A(net985),
    .B(net986),
    .C(_03814_),
    .Y(_03816_));
 sg13g2_or2_1 _09811_ (.X(_03817_),
    .B(_03816_),
    .A(net919));
 sg13g2_buf_1 fanout906 (.A(net907),
    .X(net906));
 sg13g2_a21oi_1 _09813_ (.A1(_03805_),
    .A2(_03810_),
    .Y(_03819_),
    .B1(_03817_));
 sg13g2_buf_1 fanout905 (.A(net906),
    .X(net905));
 sg13g2_buf_2 fanout904 (.A(net906),
    .X(net904));
 sg13g2_buf_1 fanout903 (.A(_04429_),
    .X(net903));
 sg13g2_buf_2 fanout902 (.A(net903),
    .X(net902));
 sg13g2_and3_1 _09818_ (.X(_03824_),
    .A(net1),
    .B(net12),
    .C(net1248));
 sg13g2_buf_2 fanout901 (.A(net902),
    .X(net901));
 sg13g2_and3_2 _09820_ (.X(_03826_),
    .A(net1255),
    .B(_02561_),
    .C(_03824_));
 sg13g2_buf_1 fanout900 (.A(net903),
    .X(net900));
 sg13g2_nor3_1 _09822_ (.A(net1249),
    .B(net986),
    .C(net1036),
    .Y(_03828_));
 sg13g2_nand2_1 _09823_ (.Y(_03829_),
    .A(net1),
    .B(net12));
 sg13g2_nor3_1 _09824_ (.A(net985),
    .B(_03829_),
    .C(_03799_),
    .Y(_03830_));
 sg13g2_nor4_2 _09825_ (.A(net919),
    .B(_03826_),
    .C(_03828_),
    .Y(_03831_),
    .D(_03830_));
 sg13g2_buf_2 fanout899 (.A(net903),
    .X(net899));
 sg13g2_buf_1 fanout898 (.A(_04436_),
    .X(net898));
 sg13g2_buf_2 fanout897 (.A(_04436_),
    .X(net897));
 sg13g2_buf_2 fanout896 (.A(_04488_),
    .X(net896));
 sg13g2_nand2_1 _09830_ (.Y(_03836_),
    .A(net1251),
    .B(net1254));
 sg13g2_a22oi_1 _09831_ (.Y(_03837_),
    .B1(_03814_),
    .B2(net985),
    .A2(_03836_),
    .A1(net986));
 sg13g2_buf_2 fanout895 (.A(_04827_),
    .X(net895));
 sg13g2_nor3_1 _09833_ (.A(net99),
    .B(net923),
    .C(_03837_),
    .Y(_03839_));
 sg13g2_buf_1 fanout894 (.A(_06778_),
    .X(net894));
 sg13g2_and2_1 _09835_ (.A(net30),
    .B(net99),
    .X(_03841_));
 sg13g2_a22oi_1 _09836_ (.Y(_03842_),
    .B1(_03841_),
    .B2(net911),
    .A2(_03839_),
    .A1(net1375));
 sg13g2_a21oi_1 _09837_ (.A1(_03448_),
    .A2(net911),
    .Y(_03843_),
    .B1(_03842_));
 sg13g2_buf_1 fanout893 (.A(net894),
    .X(net893));
 sg13g2_buf_2 fanout892 (.A(net894),
    .X(net892));
 sg13g2_buf_2 fanout891 (.A(_06778_),
    .X(net891));
 sg13g2_xnor2_1 _09841_ (.Y(_03847_),
    .A(net880),
    .B(net642));
 sg13g2_buf_2 fanout890 (.A(net891),
    .X(net890));
 sg13g2_a21oi_1 _09843_ (.A1(net1249),
    .A2(net24),
    .Y(_03849_),
    .B1(_03796_));
 sg13g2_nor2_1 _09844_ (.A(_03801_),
    .B(_03849_),
    .Y(_03850_));
 sg13g2_nor2_1 _09845_ (.A(_03817_),
    .B(_03850_),
    .Y(_03851_));
 sg13g2_nand3_1 _09846_ (.B(_02576_),
    .C(_03851_),
    .A(net1238),
    .Y(_03852_));
 sg13g2_buf_2 fanout889 (.A(net890),
    .X(net889));
 sg13g2_buf_2 fanout888 (.A(_06782_),
    .X(net888));
 sg13g2_buf_2 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_2 fanout886 (.A(net887),
    .X(net886));
 sg13g2_nor2_1 _09851_ (.A(net919),
    .B(_03816_),
    .Y(_03857_));
 sg13g2_buf_2 fanout885 (.A(net886),
    .X(net885));
 sg13g2_nand2b_1 _09853_ (.Y(_03859_),
    .B(net1243),
    .A_N(net1241));
 sg13g2_buf_2 fanout884 (.A(net886),
    .X(net884));
 sg13g2_nand2b_1 _09855_ (.Y(_03861_),
    .B(net24),
    .A_N(net1238));
 sg13g2_nor2_1 _09856_ (.A(_02576_),
    .B(_03861_),
    .Y(_03862_));
 sg13g2_a22oi_1 _09857_ (.Y(_03863_),
    .B1(_03862_),
    .B2(_03801_),
    .A2(net983),
    .A1(net1238));
 sg13g2_nand2b_1 _09858_ (.Y(_03864_),
    .B(_03863_),
    .A_N(_03806_));
 sg13g2_nor2_1 _09859_ (.A(net27),
    .B(_03801_),
    .Y(_03865_));
 sg13g2_nand3_1 _09860_ (.B(net1239),
    .C(_03865_),
    .A(net1242),
    .Y(_03866_));
 sg13g2_buf_2 fanout883 (.A(net888),
    .X(net883));
 sg13g2_buf_1 fanout882 (.A(_03819_),
    .X(net882));
 sg13g2_buf_2 fanout881 (.A(net882),
    .X(net881));
 sg13g2_nor2_1 _09864_ (.A(net986),
    .B(net1036),
    .Y(_03870_));
 sg13g2_nor2b_1 _09865_ (.A(net1242),
    .B_N(net1237),
    .Y(_03871_));
 sg13g2_a21oi_1 _09866_ (.A1(net1249),
    .A2(_03870_),
    .Y(_03872_),
    .B1(_03871_));
 sg13g2_nand2b_1 _09867_ (.Y(_03873_),
    .B(net27),
    .A_N(_03872_));
 sg13g2_nor2_1 _09868_ (.A(net1242),
    .B(_03870_),
    .Y(_03874_));
 sg13g2_o21ai_1 _09869_ (.B1(net1237),
    .Y(_03875_),
    .A1(net1239),
    .A2(_03874_));
 sg13g2_nand3_1 _09870_ (.B(_03873_),
    .C(_03875_),
    .A(_03866_),
    .Y(_03876_));
 sg13g2_and3_1 _09871_ (.X(_03877_),
    .A(_03857_),
    .B(_03864_),
    .C(_03876_));
 sg13g2_buf_2 fanout880 (.A(_03819_),
    .X(net880));
 sg13g2_buf_1 fanout879 (.A(net880),
    .X(net879));
 sg13g2_nand2_1 _09874_ (.Y(_03880_),
    .A(net849),
    .B(net635));
 sg13g2_nand2_1 _09875_ (.Y(_03881_),
    .A(net1237),
    .B(net1242));
 sg13g2_nand3_1 _09876_ (.B(_03851_),
    .C(_03881_),
    .A(net1240),
    .Y(_03882_));
 sg13g2_buf_2 fanout878 (.A(net879),
    .X(net878));
 sg13g2_buf_1 fanout877 (.A(_04055_),
    .X(net877));
 sg13g2_o21ai_1 _09879_ (.B1(net844),
    .Y(_03885_),
    .A1(_03847_),
    .A2(_03880_));
 sg13g2_a21oi_1 _09880_ (.A1(_03847_),
    .A2(net635),
    .Y(_03886_),
    .B1(net844));
 sg13g2_a21oi_1 _09881_ (.A1(net648),
    .A2(_03885_),
    .Y(_03887_),
    .B1(_03886_));
 sg13g2_buf_2 fanout876 (.A(net877),
    .X(net876));
 sg13g2_nand2_1 _09883_ (.Y(_03889_),
    .A(_03049_),
    .B(_03331_));
 sg13g2_xnor2_1 _09884_ (.Y(_03890_),
    .A(net878),
    .B(_03889_));
 sg13g2_buf_2 fanout875 (.A(net876),
    .X(net875));
 sg13g2_buf_4 fanout874 (.X(net874),
    .A(net875));
 sg13g2_and2_2 _09887_ (.A(net25),
    .B(net933),
    .X(_03893_));
 sg13g2_buf_2 fanout873 (.A(net877),
    .X(net873));
 sg13g2_a21o_2 _09889_ (.A2(net918),
    .A1(net1338),
    .B1(_03893_),
    .X(_03895_));
 sg13g2_buf_4 fanout872 (.X(net872),
    .A(net877));
 sg13g2_a21o_1 _09891_ (.A2(net918),
    .A1(net20),
    .B1(_03893_),
    .X(_03897_));
 sg13g2_buf_2 fanout871 (.A(_05453_),
    .X(net871));
 sg13g2_nor2_1 _09893_ (.A(net878),
    .B(_03897_),
    .Y(_03899_));
 sg13g2_a22oi_1 _09894_ (.Y(_03900_),
    .B1(_03899_),
    .B2(net905),
    .A2(_03895_),
    .A1(net878));
 sg13g2_a21o_1 _09895_ (.A2(_03890_),
    .A1(net904),
    .B1(_03900_),
    .X(_03901_));
 sg13g2_buf_2 fanout870 (.A(_05709_),
    .X(net870));
 sg13g2_inv_1 _09897_ (.Y(_03903_),
    .A(_03901_));
 sg13g2_buf_2 fanout869 (.A(net870),
    .X(net869));
 sg13g2_buf_2 fanout868 (.A(_05709_),
    .X(net868));
 sg13g2_buf_2 fanout867 (.A(_05810_),
    .X(net867));
 sg13g2_buf_2 fanout866 (.A(_05810_),
    .X(net866));
 sg13g2_buf_1 fanout865 (.A(_05810_),
    .X(net865));
 sg13g2_buf_1 fanout864 (.A(net865),
    .X(net864));
 sg13g2_o21ai_1 _09904_ (.B1(net1142),
    .Y(_03910_),
    .A1(net1028),
    .A2(net1014));
 sg13g2_mux2_1 _09905_ (.A0(_00162_),
    .A1(_00160_),
    .S(_03910_),
    .X(_03911_));
 sg13g2_nand3_1 _09906_ (.B(net1040),
    .C(_03911_),
    .A(net1002),
    .Y(_03912_));
 sg13g2_buf_1 fanout863 (.A(net864),
    .X(net863));
 sg13g2_buf_2 fanout862 (.A(net863),
    .X(net862));
 sg13g2_inv_1 _09909_ (.Y(_03915_),
    .A(_00174_));
 sg13g2_o21ai_1 _09910_ (.B1(_03915_),
    .Y(_03916_),
    .A1(net1026),
    .A2(net1012));
 sg13g2_inv_2 _09911_ (.Y(_03917_),
    .A(net1206));
 sg13g2_buf_2 fanout861 (.A(_07403_),
    .X(net861));
 sg13g2_buf_2 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_2 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_1 fanout858 (.A(_07403_),
    .X(net858));
 sg13g2_buf_2 fanout857 (.A(net858),
    .X(net857));
 sg13g2_buf_2 fanout856 (.A(_07427_),
    .X(net856));
 sg13g2_mux4_1 _09918_ (.S0(net970),
    .A0(_00173_),
    .A1(_00172_),
    .A2(_00175_),
    .A3(_03916_),
    .S1(net1132),
    .X(_03924_));
 sg13g2_o21ai_1 _09919_ (.B1(net1396),
    .Y(_03925_),
    .A1(net1026),
    .A2(net1012));
 sg13g2_buf_2 fanout855 (.A(net856),
    .X(net855));
 sg13g2_buf_1 fanout854 (.A(_07427_),
    .X(net854));
 sg13g2_buf_2 fanout853 (.A(_07427_),
    .X(net853));
 sg13g2_buf_1 fanout852 (.A(_03852_),
    .X(net852));
 sg13g2_buf_2 fanout851 (.A(net852),
    .X(net851));
 sg13g2_mux4_1 _09925_ (.S0(net1125),
    .A0(_00168_),
    .A1(_00170_),
    .A2(_00169_),
    .A3(_00171_),
    .S1(net1205),
    .X(_03931_));
 sg13g2_nor2_1 _09926_ (.A(net1106),
    .B(_03931_),
    .Y(_03932_));
 sg13g2_nor2_1 _09927_ (.A(_03925_),
    .B(_03932_),
    .Y(_03933_));
 sg13g2_inv_1 _09928_ (.Y(_03934_),
    .A(_00164_));
 sg13g2_nor2b_2 _09929_ (.A(net1221),
    .B_N(net1110),
    .Y(_03935_));
 sg13g2_buf_2 fanout850 (.A(net851),
    .X(net850));
 sg13g2_nand2_1 _09931_ (.Y(_03937_),
    .A(net1106),
    .B(_00165_));
 sg13g2_buf_1 fanout849 (.A(net852),
    .X(net849));
 sg13g2_buf_2 fanout848 (.A(net852),
    .X(net848));
 sg13g2_buf_1 fanout847 (.A(_03882_),
    .X(net847));
 sg13g2_buf_2 fanout846 (.A(net847),
    .X(net846));
 sg13g2_buf_2 fanout845 (.A(net846),
    .X(net845));
 sg13g2_a221oi_1 _09937_ (.B2(net1208),
    .C1(net1132),
    .B1(_03937_),
    .A1(_03934_),
    .Y(_03943_),
    .A2(_03935_));
 sg13g2_buf_1 fanout844 (.A(_03882_),
    .X(net844));
 sg13g2_buf_1 fanout843 (.A(net844),
    .X(net843));
 sg13g2_buf_1 fanout842 (.A(net843),
    .X(net842));
 sg13g2_mux2_1 _09941_ (.A0(_00166_),
    .A1(_00167_),
    .S(net1213),
    .X(_03947_));
 sg13g2_nand3_1 _09942_ (.B(net1109),
    .C(_03947_),
    .A(net1133),
    .Y(_03948_));
 sg13g2_nand2b_1 _09943_ (.Y(_03949_),
    .B(_03948_),
    .A_N(_03943_));
 sg13g2_buf_2 fanout841 (.A(net843),
    .X(net841));
 sg13g2_o21ai_1 _09945_ (.B1(net996),
    .Y(_03951_),
    .A1(net1035),
    .A2(net1021));
 sg13g2_and2_1 _09946_ (.A(net992),
    .B(_03931_),
    .X(_03952_));
 sg13g2_buf_1 fanout840 (.A(_05785_),
    .X(net840));
 sg13g2_buf_1 fanout839 (.A(net840),
    .X(net839));
 sg13g2_nand2_1 _09949_ (.Y(_03955_),
    .A(net1142),
    .B(_00163_));
 sg13g2_buf_2 fanout838 (.A(net840),
    .X(net838));
 sg13g2_buf_1 fanout837 (.A(net840),
    .X(net837));
 sg13g2_nand2b_1 _09952_ (.Y(_03958_),
    .B(_00161_),
    .A_N(net1142));
 sg13g2_buf_2 fanout836 (.A(net837),
    .X(net836));
 sg13g2_buf_2 fanout835 (.A(net837),
    .X(net835));
 sg13g2_a22oi_1 _09955_ (.Y(_03961_),
    .B1(net1396),
    .B2(net1004),
    .A2(_03958_),
    .A1(_03955_));
 sg13g2_or3_1 _09956_ (.A(_03951_),
    .B(_03952_),
    .C(_03961_),
    .X(_03962_));
 sg13g2_a221oi_1 _09957_ (.B2(net1002),
    .C1(_03962_),
    .B1(_03949_),
    .A1(_03924_),
    .Y(_03963_),
    .A2(_03933_));
 sg13g2_and2_1 _09958_ (.A(net1106),
    .B(net1396),
    .X(_03964_));
 sg13g2_buf_2 fanout834 (.A(_05804_),
    .X(net834));
 sg13g2_buf_2 fanout833 (.A(net834),
    .X(net833));
 sg13g2_buf_2 fanout832 (.A(_05804_),
    .X(net832));
 sg13g2_buf_2 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_2 fanout830 (.A(net832),
    .X(net830));
 sg13g2_mux4_1 _09964_ (.S0(net1126),
    .A0(_00188_),
    .A1(_00190_),
    .A2(_00189_),
    .A3(_00191_),
    .S1(net1205),
    .X(_03970_));
 sg13g2_buf_2 fanout829 (.A(net98),
    .X(net829));
 sg13g2_a21oi_1 _09966_ (.A1(net969),
    .A2(_03970_),
    .Y(_03972_),
    .B1(net945));
 sg13g2_nor2b_1 _09967_ (.A(net1396),
    .B_N(net1106),
    .Y(_03973_));
 sg13g2_buf_2 fanout828 (.A(net829),
    .X(net828));
 sg13g2_buf_2 fanout827 (.A(net828),
    .X(net827));
 sg13g2_buf_1 fanout826 (.A(_05814_),
    .X(net826));
 sg13g2_buf_1 fanout825 (.A(net826),
    .X(net825));
 sg13g2_mux4_1 _09972_ (.S0(net1126),
    .A0(_00180_),
    .A1(_00182_),
    .A2(_00181_),
    .A3(_00183_),
    .S1(net1205),
    .X(_03978_));
 sg13g2_mux4_1 _09973_ (.S0(net1127),
    .A0(_00176_),
    .A1(_00178_),
    .A2(_00177_),
    .A3(_00179_),
    .S1(net1205),
    .X(_03979_));
 sg13g2_nor2_1 _09974_ (.A(net1106),
    .B(net1396),
    .Y(_03980_));
 sg13g2_buf_2 fanout824 (.A(net825),
    .X(net824));
 sg13g2_buf_2 fanout823 (.A(net826),
    .X(net823));
 sg13g2_buf_1 fanout822 (.A(_05902_),
    .X(net822));
 sg13g2_buf_1 fanout821 (.A(net822),
    .X(net821));
 sg13g2_mux4_1 _09979_ (.S0(net1126),
    .A0(_00184_),
    .A1(_00186_),
    .A2(_00185_),
    .A3(_00187_),
    .S1(net1205),
    .X(_03985_));
 sg13g2_and2_1 _09980_ (.A(net992),
    .B(_03985_),
    .X(_03986_));
 sg13g2_a221oi_1 _09981_ (.B2(net963),
    .C1(_03986_),
    .B1(_03979_),
    .A1(net966),
    .Y(_03987_),
    .A2(_03978_));
 sg13g2_and2_1 _09982_ (.A(_03972_),
    .B(_03987_),
    .X(_03988_));
 sg13g2_a21oi_2 _09983_ (.B1(_03988_),
    .Y(_03989_),
    .A2(_03963_),
    .A1(_03912_));
 sg13g2_buf_2 fanout820 (.A(net822),
    .X(net820));
 sg13g2_buf_1 fanout819 (.A(_05902_),
    .X(net819));
 sg13g2_buf_1 fanout818 (.A(net819),
    .X(net818));
 sg13g2_buf_1 fanout817 (.A(net818),
    .X(net817));
 sg13g2_buf_2 fanout816 (.A(net818),
    .X(net816));
 sg13g2_or2_1 _09989_ (.X(_03995_),
    .B(_00256_),
    .A(net1151));
 sg13g2_buf_2 fanout815 (.A(_06020_),
    .X(net815));
 sg13g2_nor2b_1 _09991_ (.A(_00258_),
    .B_N(net1151),
    .Y(_03997_));
 sg13g2_o21ai_1 _09992_ (.B1(_03997_),
    .Y(_03998_),
    .A1(net1027),
    .A2(net1013));
 sg13g2_buf_2 fanout814 (.A(_06020_),
    .X(net814));
 sg13g2_a21o_1 _09994_ (.A2(_03998_),
    .A1(_03995_),
    .B1(net1216),
    .X(_04000_));
 sg13g2_buf_2 fanout813 (.A(_07434_),
    .X(net813));
 sg13g2_buf_2 fanout812 (.A(net813),
    .X(net812));
 sg13g2_buf_2 fanout811 (.A(net813),
    .X(net811));
 sg13g2_mux2_1 _09998_ (.A0(_00257_),
    .A1(_00259_),
    .S(net1151),
    .X(_04004_));
 sg13g2_o21ai_1 _09999_ (.B1(net964),
    .Y(_04005_),
    .A1(net974),
    .A2(_04004_));
 sg13g2_nor3_1 _10000_ (.A(_00256_),
    .B(net1030),
    .C(net1016),
    .Y(_04006_));
 sg13g2_a21oi_1 _10001_ (.A1(net926),
    .A2(_04005_),
    .Y(_04007_),
    .B1(_04006_));
 sg13g2_buf_2 fanout810 (.A(net811),
    .X(net810));
 sg13g2_a21oi_2 _10003_ (.B1(net1392),
    .Y(_04009_),
    .A2(_03743_),
    .A1(net963));
 sg13g2_buf_2 fanout809 (.A(net813),
    .X(net809));
 sg13g2_mux4_1 _10005_ (.S0(net1130),
    .A0(_00260_),
    .A1(_00262_),
    .A2(_00261_),
    .A3(_00263_),
    .S1(net1207),
    .X(_04011_));
 sg13g2_nand2_1 _10006_ (.Y(_04012_),
    .A(net966),
    .B(_04011_));
 sg13g2_nand3_1 _10007_ (.B(_04009_),
    .C(_04012_),
    .A(net927),
    .Y(_04013_));
 sg13g2_o21ai_1 _10008_ (.B1(_03964_),
    .Y(_04014_),
    .A1(net1027),
    .A2(net1013));
 sg13g2_buf_2 fanout808 (.A(net809),
    .X(net808));
 sg13g2_buf_1 fanout807 (.A(net808),
    .X(net807));
 sg13g2_buf_2 fanout806 (.A(net808),
    .X(net806));
 sg13g2_buf_2 fanout805 (.A(_07564_),
    .X(net805));
 sg13g2_buf_2 fanout804 (.A(net805),
    .X(net804));
 sg13g2_mux4_1 _10014_ (.S0(net1130),
    .A0(_00268_),
    .A1(_00270_),
    .A2(_00269_),
    .A3(_00271_),
    .S1(net1207),
    .X(_04020_));
 sg13g2_inv_1 _10015_ (.Y(_04021_),
    .A(_04020_));
 sg13g2_mux4_1 _10016_ (.S0(net1151),
    .A0(_00264_),
    .A1(_00266_),
    .A2(_00265_),
    .A3(_00267_),
    .S1(net1216),
    .X(_04022_));
 sg13g2_nand2_1 _10017_ (.Y(_04023_),
    .A(net991),
    .B(_04022_));
 sg13g2_o21ai_1 _10018_ (.B1(_04023_),
    .Y(_04024_),
    .A1(_04014_),
    .A2(_04021_));
 sg13g2_a22oi_1 _10019_ (.Y(_04025_),
    .B1(_04013_),
    .B2(_04024_),
    .A2(_04007_),
    .A1(_04000_));
 sg13g2_or2_1 _10020_ (.X(_04026_),
    .B(_00272_),
    .A(net1130));
 sg13g2_nor2b_1 _10021_ (.A(_00274_),
    .B_N(net1130),
    .Y(_04027_));
 sg13g2_o21ai_1 _10022_ (.B1(_04027_),
    .Y(_04028_),
    .A1(net1026),
    .A2(net1012));
 sg13g2_a21o_1 _10023_ (.A2(_04028_),
    .A1(_04026_),
    .B1(net1207),
    .X(_04029_));
 sg13g2_mux2_1 _10024_ (.A0(_00273_),
    .A1(_00275_),
    .S(net1130),
    .X(_04030_));
 sg13g2_o21ai_1 _10025_ (.B1(net963),
    .Y(_04031_),
    .A1(net971),
    .A2(_04030_));
 sg13g2_nor3_1 _10026_ (.A(_00272_),
    .B(net1026),
    .C(net1012),
    .Y(_04032_));
 sg13g2_a21oi_1 _10027_ (.A1(net927),
    .A2(_04031_),
    .Y(_04033_),
    .B1(_04032_));
 sg13g2_mux4_1 _10028_ (.S0(net1151),
    .A0(_00276_),
    .A1(_00278_),
    .A2(_00277_),
    .A3(_00279_),
    .S1(net1216),
    .X(_04034_));
 sg13g2_buf_1 fanout803 (.A(_07843_),
    .X(net803));
 sg13g2_mux4_1 _10030_ (.S0(net1133),
    .A0(_00284_),
    .A1(_00286_),
    .A2(_00285_),
    .A3(_00287_),
    .S1(net1209),
    .X(_04036_));
 sg13g2_and2_1 _10031_ (.A(net969),
    .B(_04036_),
    .X(_04037_));
 sg13g2_nand2_1 _10032_ (.Y(_04038_),
    .A(net1130),
    .B(_00282_));
 sg13g2_nand2b_1 _10033_ (.Y(_04039_),
    .B(_00280_),
    .A_N(net1133));
 sg13g2_buf_1 fanout802 (.A(net803),
    .X(net802));
 sg13g2_buf_1 fanout801 (.A(net802),
    .X(net801));
 sg13g2_a22oi_1 _10036_ (.Y(_04042_),
    .B1(net1003),
    .B2(net1001),
    .A2(_04039_),
    .A1(_04038_));
 sg13g2_nand2_1 _10037_ (.Y(_04043_),
    .A(net1130),
    .B(_00283_));
 sg13g2_nand2b_1 _10038_ (.Y(_04044_),
    .B(_00281_),
    .A_N(net1133));
 sg13g2_nand3b_1 _10039_ (.B(net1398),
    .C(net1217),
    .Y(_04045_),
    .A_N(net1110));
 sg13g2_buf_2 fanout800 (.A(net802),
    .X(net800));
 sg13g2_a21oi_1 _10041_ (.A1(_04043_),
    .A2(_04044_),
    .Y(_04047_),
    .B1(_04045_));
 sg13g2_or4_1 _10042_ (.A(net945),
    .B(_04037_),
    .C(_04042_),
    .D(_04047_),
    .X(_04048_));
 sg13g2_a221oi_1 _10043_ (.B2(net967),
    .C1(_04048_),
    .B1(_04034_),
    .A1(_04029_),
    .Y(_04049_),
    .A2(_04033_));
 sg13g2_or2_1 _10044_ (.X(_04050_),
    .B(_04049_),
    .A(_04025_));
 sg13g2_buf_1 fanout799 (.A(net802),
    .X(net799));
 sg13g2_a21oi_2 _10046_ (.B1(_03893_),
    .Y(_04052_),
    .A2(net918),
    .A1(net1339));
 sg13g2_a21o_1 _10047_ (.A2(net918),
    .A1(net1259),
    .B1(_03893_),
    .X(_04053_));
 sg13g2_buf_1 fanout798 (.A(net799),
    .X(net798));
 sg13g2_a21o_1 _10049_ (.A2(_03810_),
    .A1(_03805_),
    .B1(_03817_),
    .X(_04055_));
 sg13g2_buf_2 fanout797 (.A(net799),
    .X(net797));
 sg13g2_buf_2 fanout796 (.A(net799),
    .X(net796));
 sg13g2_mux2_1 _10052_ (.A0(_04052_),
    .A1(_04053_),
    .S(net872),
    .X(_04058_));
 sg13g2_xnor2_1 _10053_ (.Y(_04059_),
    .A(_03264_),
    .B(net879));
 sg13g2_mux2_1 _10054_ (.A0(_04058_),
    .A1(_04059_),
    .S(net905),
    .X(_04060_));
 sg13g2_buf_2 fanout795 (.A(net803),
    .X(net795));
 sg13g2_nand2_1 _10056_ (.Y(_04062_),
    .A(_04050_),
    .B(_04060_));
 sg13g2_or2_1 _10057_ (.X(_04063_),
    .B(_00224_),
    .A(net1128));
 sg13g2_nor2b_1 _10058_ (.A(_00226_),
    .B_N(net1129),
    .Y(_04064_));
 sg13g2_o21ai_1 _10059_ (.B1(_04064_),
    .Y(_04065_),
    .A1(net1025),
    .A2(net1011));
 sg13g2_a21o_1 _10060_ (.A2(_04065_),
    .A1(_04063_),
    .B1(net1207),
    .X(_04066_));
 sg13g2_mux2_1 _10061_ (.A0(_00225_),
    .A1(_00227_),
    .S(net1124),
    .X(_04067_));
 sg13g2_o21ai_1 _10062_ (.B1(net963),
    .Y(_04068_),
    .A1(net970),
    .A2(_04067_));
 sg13g2_nor3_1 _10063_ (.A(_00224_),
    .B(net1025),
    .C(net1011),
    .Y(_04069_));
 sg13g2_a21oi_1 _10064_ (.A1(net926),
    .A2(_04068_),
    .Y(_04070_),
    .B1(_04069_));
 sg13g2_mux4_1 _10065_ (.S0(net1124),
    .A0(_00228_),
    .A1(_00230_),
    .A2(_00229_),
    .A3(_00231_),
    .S1(net1206),
    .X(_04071_));
 sg13g2_nand2_1 _10066_ (.Y(_04072_),
    .A(net966),
    .B(_04071_));
 sg13g2_nand3_1 _10067_ (.B(_04009_),
    .C(_04072_),
    .A(net926),
    .Y(_04073_));
 sg13g2_mux4_1 _10068_ (.S0(net1124),
    .A0(_00236_),
    .A1(_00238_),
    .A2(_00237_),
    .A3(_00239_),
    .S1(net1206),
    .X(_04074_));
 sg13g2_inv_1 _10069_ (.Y(_04075_),
    .A(_04074_));
 sg13g2_mux4_1 _10070_ (.S0(net1124),
    .A0(_00232_),
    .A1(_00234_),
    .A2(_00233_),
    .A3(_00235_),
    .S1(net1206),
    .X(_04076_));
 sg13g2_nand2_1 _10071_ (.Y(_04077_),
    .A(net992),
    .B(_04076_));
 sg13g2_o21ai_1 _10072_ (.B1(_04077_),
    .Y(_04078_),
    .A1(_04014_),
    .A2(_04075_));
 sg13g2_a22oi_1 _10073_ (.Y(_04079_),
    .B1(_04073_),
    .B2(_04078_),
    .A2(_04070_),
    .A1(_04066_));
 sg13g2_or2_1 _10074_ (.X(_04080_),
    .B(_00240_),
    .A(net1124));
 sg13g2_nor2b_1 _10075_ (.A(_00242_),
    .B_N(net1124),
    .Y(_04081_));
 sg13g2_o21ai_1 _10076_ (.B1(_04081_),
    .Y(_04082_),
    .A1(net1025),
    .A2(net1011));
 sg13g2_a21o_1 _10077_ (.A2(_04082_),
    .A1(_04080_),
    .B1(net1206),
    .X(_04083_));
 sg13g2_mux2_1 _10078_ (.A0(_00241_),
    .A1(_00243_),
    .S(net1124),
    .X(_04084_));
 sg13g2_o21ai_1 _10079_ (.B1(net963),
    .Y(_04085_),
    .A1(net970),
    .A2(_04084_));
 sg13g2_nor3_1 _10080_ (.A(_00240_),
    .B(net1025),
    .C(net1011),
    .Y(_04086_));
 sg13g2_a21oi_1 _10081_ (.A1(net926),
    .A2(_04085_),
    .Y(_04087_),
    .B1(_04086_));
 sg13g2_mux4_1 _10082_ (.S0(net1124),
    .A0(_00244_),
    .A1(_00246_),
    .A2(_00245_),
    .A3(_00247_),
    .S1(net1206),
    .X(_04088_));
 sg13g2_buf_2 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_2 fanout793 (.A(net803),
    .X(net793));
 sg13g2_mux4_1 _10085_ (.S0(net1126),
    .A0(_00252_),
    .A1(_00254_),
    .A2(_00253_),
    .A3(_00255_),
    .S1(net1205),
    .X(_04091_));
 sg13g2_and2_1 _10086_ (.A(net969),
    .B(_04091_),
    .X(_04092_));
 sg13g2_nand2_1 _10087_ (.Y(_04093_),
    .A(net1125),
    .B(_00250_));
 sg13g2_nand2b_1 _10088_ (.Y(_04094_),
    .B(_00248_),
    .A_N(net1125));
 sg13g2_a22oi_1 _10089_ (.Y(_04095_),
    .B1(net1002),
    .B2(net1001),
    .A2(_04094_),
    .A1(_04093_));
 sg13g2_nand2_1 _10090_ (.Y(_04096_),
    .A(net1127),
    .B(_00251_));
 sg13g2_nand2b_1 _10091_ (.Y(_04097_),
    .B(_00249_),
    .A_N(net1125));
 sg13g2_a21oi_1 _10092_ (.A1(_04096_),
    .A2(_04097_),
    .Y(_04098_),
    .B1(_04045_));
 sg13g2_or4_1 _10093_ (.A(net945),
    .B(_04092_),
    .C(_04095_),
    .D(_04098_),
    .X(_04099_));
 sg13g2_a221oi_1 _10094_ (.B2(net966),
    .C1(_04099_),
    .B1(_04088_),
    .A1(_04083_),
    .Y(_04100_),
    .A2(_04087_));
 sg13g2_nor2_1 _10095_ (.A(_04079_),
    .B(_04100_),
    .Y(_04101_));
 sg13g2_buf_2 fanout792 (.A(net803),
    .X(net792));
 sg13g2_inv_1 _10097_ (.Y(_04103_),
    .A(net18));
 sg13g2_o21ai_1 _10098_ (.B1(net25),
    .Y(_04104_),
    .A1(net1033),
    .A2(net1019));
 sg13g2_buf_1 fanout791 (.A(_07932_),
    .X(net791));
 sg13g2_o21ai_1 _10100_ (.B1(_04104_),
    .Y(_04106_),
    .A1(_04103_),
    .A2(net931));
 sg13g2_buf_1 fanout790 (.A(net791),
    .X(net790));
 sg13g2_nor2_1 _10102_ (.A(net904),
    .B(_04106_),
    .Y(_04108_));
 sg13g2_a21oi_1 _10103_ (.A1(_03296_),
    .A2(net905),
    .Y(_04109_),
    .B1(_04108_));
 sg13g2_xnor2_1 _10104_ (.Y(_04110_),
    .A(net872),
    .B(_04109_));
 sg13g2_nand2b_1 _10105_ (.Y(_04111_),
    .B(_04110_),
    .A_N(net633));
 sg13g2_nor2b_1 _10106_ (.A(_04110_),
    .B_N(net633),
    .Y(_04112_));
 sg13g2_a21oi_2 _10107_ (.B1(_04112_),
    .Y(_04113_),
    .A2(_04111_),
    .A1(_04062_));
 sg13g2_buf_2 fanout789 (.A(net791),
    .X(net789));
 sg13g2_o21ai_1 _10109_ (.B1(net966),
    .Y(_04115_),
    .A1(net1026),
    .A2(net1012));
 sg13g2_buf_2 fanout788 (.A(net791),
    .X(net788));
 sg13g2_buf_1 fanout787 (.A(net788),
    .X(net787));
 sg13g2_inv_1 _10112_ (.Y(_04118_),
    .A(_00198_));
 sg13g2_o21ai_1 _10113_ (.B1(_04118_),
    .Y(_04119_),
    .A1(net1030),
    .A2(net1016));
 sg13g2_mux4_1 _10114_ (.S0(net974),
    .A0(_00197_),
    .A1(_00196_),
    .A2(_00199_),
    .A3(_04119_),
    .S1(net1150),
    .X(_04120_));
 sg13g2_nand2b_1 _10115_ (.Y(_04121_),
    .B(_04120_),
    .A_N(_04115_));
 sg13g2_or2_1 _10116_ (.X(_04122_),
    .B(_00192_),
    .A(net1153));
 sg13g2_buf_2 fanout786 (.A(net788),
    .X(net786));
 sg13g2_nor2b_1 _10118_ (.A(_00194_),
    .B_N(net1153),
    .Y(_04124_));
 sg13g2_o21ai_1 _10119_ (.B1(_04124_),
    .Y(_04125_),
    .A1(net1030),
    .A2(net1016));
 sg13g2_a21o_1 _10120_ (.A2(_04125_),
    .A1(_04122_),
    .B1(net1217),
    .X(_04126_));
 sg13g2_buf_2 fanout785 (.A(net791),
    .X(net785));
 sg13g2_buf_2 fanout784 (.A(net785),
    .X(net784));
 sg13g2_buf_2 fanout783 (.A(net784),
    .X(net783));
 sg13g2_buf_2 fanout782 (.A(_08006_),
    .X(net782));
 sg13g2_buf_2 fanout781 (.A(net782),
    .X(net781));
 sg13g2_mux2_1 _10126_ (.A0(_00193_),
    .A1(_00195_),
    .S(net1151),
    .X(_04132_));
 sg13g2_o21ai_1 _10127_ (.B1(net964),
    .Y(_04133_),
    .A1(net974),
    .A2(_04132_));
 sg13g2_nor3_1 _10128_ (.A(_00192_),
    .B(net1030),
    .C(net1016),
    .Y(_04134_));
 sg13g2_a21oi_1 _10129_ (.A1(net932),
    .A2(_04133_),
    .Y(_04135_),
    .B1(_04134_));
 sg13g2_mux4_1 _10130_ (.S0(net1151),
    .A0(_00204_),
    .A1(_00206_),
    .A2(_00205_),
    .A3(_00207_),
    .S1(net1216),
    .X(_04136_));
 sg13g2_inv_1 _10131_ (.Y(_04137_),
    .A(_04136_));
 sg13g2_mux4_1 _10132_ (.S0(net1151),
    .A0(_00200_),
    .A1(_00202_),
    .A2(_00201_),
    .A3(_00203_),
    .S1(net1216),
    .X(_04138_));
 sg13g2_nand2_1 _10133_ (.Y(_04139_),
    .A(net991),
    .B(_04138_));
 sg13g2_o21ai_1 _10134_ (.B1(_04139_),
    .Y(_04140_),
    .A1(_04014_),
    .A2(_04137_));
 sg13g2_nand2_2 _10135_ (.Y(_04141_),
    .A(net931),
    .B(_04009_));
 sg13g2_a22oi_1 _10136_ (.Y(_04142_),
    .B1(_04140_),
    .B2(_04141_),
    .A2(_04135_),
    .A1(_04126_));
 sg13g2_nand2_1 _10137_ (.Y(_04143_),
    .A(net1107),
    .B(net1397));
 sg13g2_nor2_1 _10138_ (.A(net920),
    .B(_04143_),
    .Y(_04144_));
 sg13g2_buf_2 fanout780 (.A(net782),
    .X(net780));
 sg13g2_inv_1 _10140_ (.Y(_04146_),
    .A(_00222_));
 sg13g2_o21ai_1 _10141_ (.B1(_04146_),
    .Y(_04147_),
    .A1(net1025),
    .A2(net1011));
 sg13g2_mux4_1 _10142_ (.S0(net970),
    .A0(_00221_),
    .A1(_00220_),
    .A2(_00223_),
    .A3(_04147_),
    .S1(net1126),
    .X(_04148_));
 sg13g2_or2_1 _10143_ (.X(_04149_),
    .B(_00208_),
    .A(net1125));
 sg13g2_nor2b_1 _10144_ (.A(_00210_),
    .B_N(net1125),
    .Y(_04150_));
 sg13g2_o21ai_1 _10145_ (.B1(_04150_),
    .Y(_04151_),
    .A1(net1026),
    .A2(net1012));
 sg13g2_a21o_1 _10146_ (.A2(_04151_),
    .A1(_04149_),
    .B1(net1210),
    .X(_04152_));
 sg13g2_buf_1 fanout779 (.A(net780),
    .X(net779));
 sg13g2_buf_2 fanout778 (.A(net780),
    .X(net778));
 sg13g2_mux2_1 _10149_ (.A0(_00209_),
    .A1(_00211_),
    .S(net1127),
    .X(_04155_));
 sg13g2_o21ai_1 _10150_ (.B1(net963),
    .Y(_04156_),
    .A1(net970),
    .A2(_04155_));
 sg13g2_nor3_1 _10151_ (.A(_00208_),
    .B(net1025),
    .C(net1011),
    .Y(_04157_));
 sg13g2_a21oi_1 _10152_ (.A1(net926),
    .A2(_04156_),
    .Y(_04158_),
    .B1(_04157_));
 sg13g2_buf_2 fanout777 (.A(_08006_),
    .X(net777));
 sg13g2_mux4_1 _10154_ (.S0(net1126),
    .A0(_00216_),
    .A1(_00218_),
    .A2(_00217_),
    .A3(_00219_),
    .S1(net1205),
    .X(_04160_));
 sg13g2_nand2_1 _10155_ (.Y(_04161_),
    .A(net992),
    .B(_04160_));
 sg13g2_mux4_1 _10156_ (.S0(net1126),
    .A0(_00212_),
    .A1(_00214_),
    .A2(_00213_),
    .A3(_00215_),
    .S1(net1205),
    .X(_04162_));
 sg13g2_nand2_1 _10157_ (.Y(_04163_),
    .A(net966),
    .B(_04162_));
 sg13g2_nand4_1 _10158_ (.B(net926),
    .C(_04161_),
    .A(net1392),
    .Y(_04164_),
    .D(_04163_));
 sg13g2_a221oi_1 _10159_ (.B2(_04158_),
    .C1(_04164_),
    .B1(_04152_),
    .A1(_04144_),
    .Y(_04165_),
    .A2(_04148_));
 sg13g2_a21oi_1 _10160_ (.A1(_04121_),
    .A2(_04142_),
    .Y(_04166_),
    .B1(_04165_));
 sg13g2_buf_2 fanout776 (.A(net777),
    .X(net776));
 sg13g2_inv_1 _10162_ (.Y(_04168_),
    .A(net19));
 sg13g2_o21ai_1 _10163_ (.B1(_04104_),
    .Y(_04169_),
    .A1(_04168_),
    .A2(net931));
 sg13g2_buf_1 fanout775 (.A(net776),
    .X(net775));
 sg13g2_nor2_1 _10165_ (.A(net904),
    .B(_04169_),
    .Y(_04171_));
 sg13g2_a21oi_1 _10166_ (.A1(_03314_),
    .A2(net905),
    .Y(_04172_),
    .B1(_04171_));
 sg13g2_xnor2_1 _10167_ (.Y(_04173_),
    .A(net879),
    .B(_04172_));
 sg13g2_buf_2 fanout774 (.A(net776),
    .X(net774));
 sg13g2_nor2_1 _10169_ (.A(net631),
    .B(_04173_),
    .Y(_04175_));
 sg13g2_or2_1 _10170_ (.X(_04176_),
    .B(_04175_),
    .A(_03901_));
 sg13g2_a21o_2 _10171_ (.A2(_03963_),
    .A1(_03912_),
    .B1(_03988_),
    .X(_04177_));
 sg13g2_buf_2 fanout773 (.A(_08018_),
    .X(net773));
 sg13g2_nand2_1 _10173_ (.Y(_04179_),
    .A(net631),
    .B(_04173_));
 sg13g2_a21o_1 _10174_ (.A2(_04177_),
    .A1(_03901_),
    .B1(_04179_),
    .X(_04180_));
 sg13g2_o21ai_1 _10175_ (.B1(_04180_),
    .Y(_04181_),
    .A1(_04113_),
    .A2(_04176_));
 sg13g2_nor3_1 _10176_ (.A(_04177_),
    .B(_04113_),
    .C(_04175_),
    .Y(_04182_));
 sg13g2_a22oi_1 _10177_ (.Y(_04183_),
    .B1(_04181_),
    .B2(_04182_),
    .A2(_03989_),
    .A1(_03903_));
 sg13g2_buf_2 fanout772 (.A(net773),
    .X(net772));
 sg13g2_buf_1 fanout771 (.A(_08052_),
    .X(net771));
 sg13g2_inv_1 _10180_ (.Y(_04186_),
    .A(net22));
 sg13g2_o21ai_1 _10181_ (.B1(_04104_),
    .Y(_04187_),
    .A1(_04186_),
    .A2(net933));
 sg13g2_buf_2 fanout770 (.A(net771),
    .X(net770));
 sg13g2_nor2_1 _10183_ (.A(net906),
    .B(_04187_),
    .Y(_04189_));
 sg13g2_a21oi_1 _10184_ (.A1(_03376_),
    .A2(net906),
    .Y(_04190_),
    .B1(_04189_));
 sg13g2_xnor2_1 _10185_ (.Y(_04191_),
    .A(net872),
    .B(_04190_));
 sg13g2_or2_1 _10186_ (.X(_04192_),
    .B(_00096_),
    .A(net1156));
 sg13g2_buf_2 fanout769 (.A(net771),
    .X(net769));
 sg13g2_nor2b_1 _10188_ (.A(_00098_),
    .B_N(net1156),
    .Y(_04194_));
 sg13g2_o21ai_1 _10189_ (.B1(_04194_),
    .Y(_04195_),
    .A1(net1032),
    .A2(net1018));
 sg13g2_a21o_1 _10190_ (.A2(_04195_),
    .A1(_04192_),
    .B1(net1219),
    .X(_04196_));
 sg13g2_buf_2 fanout768 (.A(net769),
    .X(net768));
 sg13g2_mux2_1 _10192_ (.A0(_00097_),
    .A1(_00099_),
    .S(net1156),
    .X(_04198_));
 sg13g2_o21ai_1 _10193_ (.B1(net964),
    .Y(_04199_),
    .A1(net975),
    .A2(_04198_));
 sg13g2_nor3_1 _10194_ (.A(_00096_),
    .B(net1032),
    .C(net1018),
    .Y(_04200_));
 sg13g2_a21oi_1 _10195_ (.A1(net931),
    .A2(_04199_),
    .Y(_04201_),
    .B1(_04200_));
 sg13g2_mux4_1 _10196_ (.S0(net1156),
    .A0(_00108_),
    .A1(_00110_),
    .A2(_00109_),
    .A3(_00111_),
    .S1(net1219),
    .X(_04202_));
 sg13g2_inv_1 _10197_ (.Y(_04203_),
    .A(_04202_));
 sg13g2_mux4_1 _10198_ (.S0(net1157),
    .A0(_00104_),
    .A1(_00106_),
    .A2(_00105_),
    .A3(_00107_),
    .S1(net1220),
    .X(_04204_));
 sg13g2_nand2_1 _10199_ (.Y(_04205_),
    .A(net991),
    .B(_04204_));
 sg13g2_o21ai_1 _10200_ (.B1(_04205_),
    .Y(_04206_),
    .A1(_04014_),
    .A2(_04203_));
 sg13g2_buf_2 fanout767 (.A(_08052_),
    .X(net767));
 sg13g2_mux4_1 _10202_ (.S0(net1157),
    .A0(_00100_),
    .A1(_00102_),
    .A2(_00101_),
    .A3(_00103_),
    .S1(net1220),
    .X(_04208_));
 sg13g2_nand2_1 _10203_ (.Y(_04209_),
    .A(net967),
    .B(_04208_));
 sg13g2_nand3_1 _10204_ (.B(_04009_),
    .C(_04209_),
    .A(net931),
    .Y(_04210_));
 sg13g2_a22oi_1 _10205_ (.Y(_04211_),
    .B1(_04206_),
    .B2(_04210_),
    .A2(_04201_),
    .A1(_04196_));
 sg13g2_buf_2 fanout766 (.A(net767),
    .X(net766));
 sg13g2_or2_1 _10207_ (.X(_04213_),
    .B(_00112_),
    .A(net1160));
 sg13g2_nor2b_1 _10208_ (.A(_00114_),
    .B_N(net1160),
    .Y(_04214_));
 sg13g2_o21ai_1 _10209_ (.B1(_04214_),
    .Y(_04215_),
    .A1(net1031),
    .A2(net1017));
 sg13g2_a21o_1 _10210_ (.A2(_04215_),
    .A1(_04213_),
    .B1(net1222),
    .X(_04216_));
 sg13g2_buf_2 fanout765 (.A(_08059_),
    .X(net765));
 sg13g2_buf_2 fanout764 (.A(_08095_),
    .X(net764));
 sg13g2_mux2_1 _10213_ (.A0(_00113_),
    .A1(_00115_),
    .S(net1155),
    .X(_04219_));
 sg13g2_o21ai_1 _10214_ (.B1(net964),
    .Y(_04220_),
    .A1(net974),
    .A2(_04219_));
 sg13g2_nor3_1 _10215_ (.A(_00112_),
    .B(net1031),
    .C(net1017),
    .Y(_04221_));
 sg13g2_a21oi_1 _10216_ (.A1(net932),
    .A2(_04220_),
    .Y(_04222_),
    .B1(_04221_));
 sg13g2_mux4_1 _10217_ (.S0(net1161),
    .A0(_00124_),
    .A1(_00126_),
    .A2(_00125_),
    .A3(_00127_),
    .S1(net1222),
    .X(_04223_));
 sg13g2_nand2_1 _10218_ (.Y(_04224_),
    .A(net1153),
    .B(_00122_));
 sg13g2_nand2b_1 _10219_ (.Y(_04225_),
    .B(_00120_),
    .A_N(net1153));
 sg13g2_a22oi_1 _10220_ (.Y(_04226_),
    .B1(net1003),
    .B2(net1001),
    .A2(_04225_),
    .A1(_04224_));
 sg13g2_nand2_1 _10221_ (.Y(_04227_),
    .A(net1153),
    .B(_00123_));
 sg13g2_nand2b_1 _10222_ (.Y(_04228_),
    .B(_00121_),
    .A_N(net1153));
 sg13g2_a21oi_1 _10223_ (.A1(_04227_),
    .A2(_04228_),
    .Y(_04229_),
    .B1(_04045_));
 sg13g2_mux4_1 _10224_ (.S0(net1153),
    .A0(_00116_),
    .A1(_00118_),
    .A2(_00117_),
    .A3(_00119_),
    .S1(net1217),
    .X(_04230_));
 sg13g2_and2_1 _10225_ (.A(net967),
    .B(_04230_),
    .X(_04231_));
 sg13g2_or4_1 _10226_ (.A(net946),
    .B(_04226_),
    .C(_04229_),
    .D(_04231_),
    .X(_04232_));
 sg13g2_a221oi_1 _10227_ (.B2(_03964_),
    .C1(_04232_),
    .B1(_04223_),
    .A1(_04216_),
    .Y(_04233_),
    .A2(_04222_));
 sg13g2_buf_2 fanout763 (.A(net764),
    .X(net763));
 sg13g2_nor2_2 _10229_ (.A(_04211_),
    .B(_04233_),
    .Y(_04235_));
 sg13g2_xnor2_1 _10230_ (.Y(_04236_),
    .A(_04191_),
    .B(_04235_));
 sg13g2_buf_2 fanout762 (.A(net764),
    .X(net762));
 sg13g2_nor2b_2 _10232_ (.A(net1225),
    .B_N(net1165),
    .Y(_04238_));
 sg13g2_buf_2 fanout761 (.A(net762),
    .X(net761));
 sg13g2_o21ai_1 _10234_ (.B1(_04238_),
    .Y(_04240_),
    .A1(net1035),
    .A2(net1021));
 sg13g2_or2_1 _10235_ (.X(_04241_),
    .B(_04240_),
    .A(_00146_));
 sg13g2_inv_1 _10236_ (.Y(_04242_),
    .A(_00144_));
 sg13g2_nor2b_1 _10237_ (.A(net1133),
    .B_N(_00145_),
    .Y(_04243_));
 sg13g2_a22oi_1 _10238_ (.Y(_04244_),
    .B1(_04243_),
    .B2(net971),
    .A2(_00147_),
    .A1(net1133));
 sg13g2_or2_2 _10239_ (.X(_04245_),
    .B(net1397),
    .A(net1109));
 sg13g2_buf_2 fanout760 (.A(_08095_),
    .X(net760));
 sg13g2_a22oi_1 _10241_ (.Y(_04247_),
    .B1(_04244_),
    .B2(_04245_),
    .A2(_03743_),
    .A1(_04242_));
 sg13g2_mux4_1 _10242_ (.S0(net1127),
    .A0(_00156_),
    .A1(_00158_),
    .A2(_00157_),
    .A3(_00159_),
    .S1(net1210),
    .X(_04248_));
 sg13g2_mux4_1 _10243_ (.S0(net1132),
    .A0(_00152_),
    .A1(_00154_),
    .A2(_00153_),
    .A3(_00155_),
    .S1(net1208),
    .X(_04249_));
 sg13g2_inv_1 _10244_ (.Y(_04250_),
    .A(net1106));
 sg13g2_buf_2 fanout759 (.A(net760),
    .X(net759));
 sg13g2_mux2_1 _10246_ (.A0(_04248_),
    .A1(_04249_),
    .S(net961),
    .X(_04252_));
 sg13g2_nand2_1 _10247_ (.Y(_04253_),
    .A(net1208),
    .B(_00151_));
 sg13g2_nand2b_1 _10248_ (.Y(_04254_),
    .B(_00150_),
    .A_N(net1208));
 sg13g2_nand3_1 _10249_ (.B(_04253_),
    .C(_04254_),
    .A(net1132),
    .Y(_04255_));
 sg13g2_inv_1 _10250_ (.Y(_04256_),
    .A(_00149_));
 sg13g2_nor2b_1 _10251_ (.A(net1132),
    .B_N(net1208),
    .Y(_04257_));
 sg13g2_nor3_1 _10252_ (.A(net1208),
    .B(net1134),
    .C(_00148_),
    .Y(_04258_));
 sg13g2_a22oi_1 _10253_ (.Y(_04259_),
    .B1(_04258_),
    .B2(_03735_),
    .A2(_04257_),
    .A1(_04256_));
 sg13g2_a21o_1 _10254_ (.A2(_04259_),
    .A1(_04255_),
    .B1(net945),
    .X(_04260_));
 sg13g2_a221oi_1 _10255_ (.B2(net1397),
    .C1(_04260_),
    .B1(_04252_),
    .A1(_04241_),
    .Y(_04261_),
    .A2(_04247_));
 sg13g2_buf_2 fanout758 (.A(net759),
    .X(net758));
 sg13g2_or2_1 _10257_ (.X(_04263_),
    .B(_04240_),
    .A(_00130_));
 sg13g2_inv_1 _10258_ (.Y(_04264_),
    .A(_00128_));
 sg13g2_nor2b_1 _10259_ (.A(net1133),
    .B_N(_00129_),
    .Y(_04265_));
 sg13g2_a22oi_1 _10260_ (.Y(_04266_),
    .B1(_04265_),
    .B2(net971),
    .A2(_00131_),
    .A1(net1133));
 sg13g2_a22oi_1 _10261_ (.Y(_04267_),
    .B1(_04266_),
    .B2(_04245_),
    .A2(_03743_),
    .A1(_04264_));
 sg13g2_mux4_1 _10262_ (.S0(net1134),
    .A0(_00136_),
    .A1(_00138_),
    .A2(_00137_),
    .A3(_00139_),
    .S1(net1209),
    .X(_04268_));
 sg13g2_nand2_1 _10263_ (.Y(_04269_),
    .A(net992),
    .B(_04268_));
 sg13g2_nand3_1 _10264_ (.B(_04009_),
    .C(_04269_),
    .A(net927),
    .Y(_04270_));
 sg13g2_mux4_1 _10265_ (.S0(net1125),
    .A0(_00132_),
    .A1(_00134_),
    .A2(_00133_),
    .A3(_00135_),
    .S1(net1210),
    .X(_04271_));
 sg13g2_nand2_1 _10266_ (.Y(_04272_),
    .A(net966),
    .B(_04271_));
 sg13g2_mux4_1 _10267_ (.S0(net1127),
    .A0(_00140_),
    .A1(_00142_),
    .A2(_00141_),
    .A3(_00143_),
    .S1(net1206),
    .X(_04273_));
 sg13g2_nand2_1 _10268_ (.Y(_04274_),
    .A(net969),
    .B(_04273_));
 sg13g2_a21oi_1 _10269_ (.A1(_04272_),
    .A2(_04274_),
    .Y(_04275_),
    .B1(net920));
 sg13g2_a22oi_1 _10270_ (.Y(_04276_),
    .B1(_04270_),
    .B2(_04275_),
    .A2(_04267_),
    .A1(_04263_));
 sg13g2_buf_2 fanout757 (.A(_08192_),
    .X(net757));
 sg13g2_or2_2 _10272_ (.X(_04278_),
    .B(_04276_),
    .A(_04261_));
 sg13g2_buf_2 fanout756 (.A(net757),
    .X(net756));
 sg13g2_inv_1 _10274_ (.Y(_04280_),
    .A(net21));
 sg13g2_o21ai_1 _10275_ (.B1(_04104_),
    .Y(_04281_),
    .A1(_04280_),
    .A2(net933));
 sg13g2_buf_2 fanout755 (.A(net756),
    .X(net755));
 sg13g2_nor2_1 _10277_ (.A(net904),
    .B(_04281_),
    .Y(_04283_));
 sg13g2_a21oi_1 _10278_ (.A1(_03359_),
    .A2(net904),
    .Y(_04284_),
    .B1(_04283_));
 sg13g2_xnor2_1 _10279_ (.Y(_04285_),
    .A(net872),
    .B(_04284_));
 sg13g2_buf_2 fanout754 (.A(net757),
    .X(net754));
 sg13g2_xnor2_1 _10281_ (.Y(_04287_),
    .A(_04278_),
    .B(_04285_));
 sg13g2_inv_1 _10282_ (.Y(_04288_),
    .A(_04287_));
 sg13g2_nand2_1 _10283_ (.Y(_04289_),
    .A(_04236_),
    .B(_04288_));
 sg13g2_nand2_1 _10284_ (.Y(_04290_),
    .A(net1243),
    .B(_03804_));
 sg13g2_nor2b_1 _10285_ (.A(_00048_),
    .B_N(net1391),
    .Y(_04291_));
 sg13g2_nand3_1 _10286_ (.B(net1391),
    .C(_00050_),
    .A(net1135),
    .Y(_04292_));
 sg13g2_o21ai_1 _10287_ (.B1(_04292_),
    .Y(_04293_),
    .A1(net1135),
    .A2(_04291_));
 sg13g2_nand2_1 _10288_ (.Y(_04294_),
    .A(net1135),
    .B(_00051_));
 sg13g2_nand2b_1 _10289_ (.Y(_04295_),
    .B(_00049_),
    .A_N(net1135));
 sg13g2_a22oi_1 _10290_ (.Y(_04296_),
    .B1(net995),
    .B2(net1004),
    .A2(_04295_),
    .A1(_04294_));
 sg13g2_a22oi_1 _10291_ (.Y(_04297_),
    .B1(_04296_),
    .B2(net920),
    .A2(_04293_),
    .A1(net1040));
 sg13g2_buf_2 fanout753 (.A(net754),
    .X(net753));
 sg13g2_buf_2 fanout752 (.A(net757),
    .X(net752));
 sg13g2_mux4_1 _10294_ (.S0(net1136),
    .A0(_00052_),
    .A1(_00054_),
    .A2(_00053_),
    .A3(_00055_),
    .S1(net1211),
    .X(_04300_));
 sg13g2_nand4_1 _10295_ (.B(net1391),
    .C(net928),
    .A(net1107),
    .Y(_04301_),
    .D(_04300_));
 sg13g2_mux4_1 _10296_ (.S0(net1136),
    .A0(_00036_),
    .A1(_00038_),
    .A2(_00037_),
    .A3(_00039_),
    .S1(net1211),
    .X(_04302_));
 sg13g2_nand3_1 _10297_ (.B(net995),
    .C(_04302_),
    .A(net1107),
    .Y(_04303_));
 sg13g2_and4_1 _10298_ (.A(net1002),
    .B(_04297_),
    .C(_04301_),
    .D(_04303_),
    .X(_04304_));
 sg13g2_inv_1 _10299_ (.Y(_04305_),
    .A(net1125));
 sg13g2_buf_2 fanout751 (.A(net752),
    .X(net751));
 sg13g2_nor2_1 _10301_ (.A(net958),
    .B(_00034_),
    .Y(_04307_));
 sg13g2_nor2_1 _10302_ (.A(net1139),
    .B(_00032_),
    .Y(_04308_));
 sg13g2_a21oi_1 _10303_ (.A1(net928),
    .A2(_04307_),
    .Y(_04309_),
    .B1(_04308_));
 sg13g2_buf_2 fanout750 (.A(net751),
    .X(net750));
 sg13g2_mux2_1 _10305_ (.A0(_00033_),
    .A1(_00035_),
    .S(net1139),
    .X(_04311_));
 sg13g2_nor2_1 _10306_ (.A(net1113),
    .B(net1393),
    .Y(_04312_));
 sg13g2_o21ai_1 _10307_ (.B1(_04312_),
    .Y(_04313_),
    .A1(net972),
    .A2(_04311_));
 sg13g2_nor3_1 _10308_ (.A(_00032_),
    .B(net1028),
    .C(net1014),
    .Y(_04314_));
 sg13g2_a21oi_1 _10309_ (.A1(net928),
    .A2(_04313_),
    .Y(_04315_),
    .B1(_04314_));
 sg13g2_o21ai_1 _10310_ (.B1(_04315_),
    .Y(_04316_),
    .A1(net1212),
    .A2(_04309_));
 sg13g2_buf_2 fanout749 (.A(net751),
    .X(net749));
 sg13g2_nor2b_1 _10312_ (.A(net1137),
    .B_N(_00060_),
    .Y(_04318_));
 sg13g2_a22oi_1 _10313_ (.Y(_04319_),
    .B1(net1007),
    .B2(_04318_),
    .A2(_00062_),
    .A1(net1137));
 sg13g2_nor2b_1 _10314_ (.A(net1138),
    .B_N(_00061_),
    .Y(_04320_));
 sg13g2_a22oi_1 _10315_ (.Y(_04321_),
    .B1(net1006),
    .B2(_04320_),
    .A2(_00063_),
    .A1(net1138));
 sg13g2_nor2b_1 _10316_ (.A(net1137),
    .B_N(_00056_),
    .Y(_04322_));
 sg13g2_a22oi_1 _10317_ (.Y(_04323_),
    .B1(net1001),
    .B2(_04322_),
    .A2(_00058_),
    .A1(net1137));
 sg13g2_nor2b_1 _10318_ (.A(net1136),
    .B_N(_00057_),
    .Y(_04324_));
 sg13g2_a22oi_1 _10319_ (.Y(_04325_),
    .B1(net1004),
    .B2(_04324_),
    .A2(_00059_),
    .A1(net1137));
 sg13g2_nor4_1 _10320_ (.A(_04319_),
    .B(_04321_),
    .C(_04323_),
    .D(_04325_),
    .Y(_04326_));
 sg13g2_or2_1 _10321_ (.X(_04327_),
    .B(_00040_),
    .A(net1139));
 sg13g2_nor2b_1 _10322_ (.A(_00042_),
    .B_N(net1136),
    .Y(_04328_));
 sg13g2_o21ai_1 _10323_ (.B1(_04328_),
    .Y(_04329_),
    .A1(net1028),
    .A2(net1014));
 sg13g2_a21o_1 _10324_ (.A2(_04329_),
    .A1(_04327_),
    .B1(net1212),
    .X(_04330_));
 sg13g2_mux2_1 _10325_ (.A0(_00041_),
    .A1(_00043_),
    .S(net1136),
    .X(_04331_));
 sg13g2_o21ai_1 _10326_ (.B1(_04312_),
    .Y(_04332_),
    .A1(net972),
    .A2(_04331_));
 sg13g2_nor3_1 _10327_ (.A(_00040_),
    .B(net1028),
    .C(net1014),
    .Y(_04333_));
 sg13g2_a21oi_1 _10328_ (.A1(net928),
    .A2(_04332_),
    .Y(_04334_),
    .B1(_04333_));
 sg13g2_nand2_1 _10329_ (.Y(_04335_),
    .A(net1137),
    .B(_00047_));
 sg13g2_nand2b_1 _10330_ (.Y(_04336_),
    .B(_00045_),
    .A_N(net1137));
 sg13g2_a22oi_1 _10331_ (.Y(_04337_),
    .B1(net1391),
    .B2(net1006),
    .A2(_04336_),
    .A1(_04335_));
 sg13g2_nand2_1 _10332_ (.Y(_04338_),
    .A(net1137),
    .B(_00046_));
 sg13g2_nand2b_1 _10333_ (.Y(_04339_),
    .B(_00044_),
    .A_N(net1138));
 sg13g2_a22oi_1 _10334_ (.Y(_04340_),
    .B1(net1391),
    .B2(net1007),
    .A2(_04339_),
    .A1(_04338_));
 sg13g2_or3_1 _10335_ (.A(_03925_),
    .B(_04337_),
    .C(_04340_),
    .X(_04341_));
 sg13g2_a221oi_1 _10336_ (.B2(_04334_),
    .C1(_04341_),
    .B1(_04330_),
    .A1(net1391),
    .Y(_04342_),
    .A2(_04326_));
 sg13g2_a21oi_1 _10337_ (.A1(_04304_),
    .A2(_04316_),
    .Y(_04343_),
    .B1(_04342_));
 sg13g2_buf_2 fanout748 (.A(_08233_),
    .X(net748));
 sg13g2_buf_2 fanout747 (.A(net748),
    .X(net747));
 sg13g2_nor2_1 _10340_ (.A(net25),
    .B(net907),
    .Y(_04346_));
 sg13g2_a21oi_2 _10341_ (.B1(_04346_),
    .Y(_04347_),
    .A2(net907),
    .A1(_03418_));
 sg13g2_xnor2_1 _10342_ (.Y(_04348_),
    .A(net630),
    .B(_04347_));
 sg13g2_o21ai_1 _10343_ (.B1(_04348_),
    .Y(_04349_),
    .A1(_03850_),
    .A2(_04290_));
 sg13g2_xnor2_1 _10344_ (.Y(_04350_),
    .A(net873),
    .B(_04349_));
 sg13g2_buf_2 fanout746 (.A(net747),
    .X(net746));
 sg13g2_xnor2_1 _10346_ (.Y(_04352_),
    .A(net880),
    .B(_04347_));
 sg13g2_nand2_1 _10347_ (.Y(_04353_),
    .A(net630),
    .B(_04352_));
 sg13g2_buf_2 fanout745 (.A(net747),
    .X(net745));
 sg13g2_or2_1 _10349_ (.X(_04355_),
    .B(_00064_),
    .A(net1219));
 sg13g2_nor2b_1 _10350_ (.A(_00065_),
    .B_N(net1219),
    .Y(_04356_));
 sg13g2_o21ai_1 _10351_ (.B1(_04356_),
    .Y(_04357_),
    .A1(net1032),
    .A2(net1018));
 sg13g2_a21o_1 _10352_ (.A2(_04357_),
    .A1(_04355_),
    .B1(net1156),
    .X(_04358_));
 sg13g2_mux2_1 _10353_ (.A0(_00066_),
    .A1(_00067_),
    .S(net1219),
    .X(_04359_));
 sg13g2_o21ai_1 _10354_ (.B1(net964),
    .Y(_04360_),
    .A1(net958),
    .A2(_04359_));
 sg13g2_nor3_1 _10355_ (.A(_00064_),
    .B(net1032),
    .C(net1018),
    .Y(_04361_));
 sg13g2_a21oi_1 _10356_ (.A1(net931),
    .A2(_04360_),
    .Y(_04362_),
    .B1(_04361_));
 sg13g2_mux4_1 _10357_ (.S0(net1157),
    .A0(_00076_),
    .A1(_00078_),
    .A2(_00077_),
    .A3(_00079_),
    .S1(net1220),
    .X(_04363_));
 sg13g2_inv_1 _10358_ (.Y(_04364_),
    .A(_04363_));
 sg13g2_mux4_1 _10359_ (.S0(net1157),
    .A0(_00068_),
    .A1(_00070_),
    .A2(_00069_),
    .A3(_00071_),
    .S1(net1220),
    .X(_04365_));
 sg13g2_nand2_1 _10360_ (.Y(_04366_),
    .A(net967),
    .B(_04365_));
 sg13g2_o21ai_1 _10361_ (.B1(_04366_),
    .Y(_04367_),
    .A1(_04364_),
    .A2(_04014_));
 sg13g2_a22oi_1 _10362_ (.Y(_04368_),
    .B1(_04141_),
    .B2(_04367_),
    .A2(_04362_),
    .A1(_04358_));
 sg13g2_inv_1 _10363_ (.Y(_04369_),
    .A(_00073_));
 sg13g2_o21ai_1 _10364_ (.B1(_04369_),
    .Y(_04370_),
    .A1(net1032),
    .A2(net1018));
 sg13g2_mux4_1 _10365_ (.S0(net1157),
    .A0(_00072_),
    .A1(_00074_),
    .A2(_04370_),
    .A3(_00075_),
    .S1(net1220),
    .X(_04371_));
 sg13g2_nand3_1 _10366_ (.B(_04371_),
    .C(net991),
    .A(net931),
    .Y(_04372_));
 sg13g2_nor2b_1 _10367_ (.A(_00089_),
    .B_N(net1221),
    .Y(_04373_));
 sg13g2_o21ai_1 _10368_ (.B1(_04373_),
    .Y(_04374_),
    .A1(net1032),
    .A2(net1018));
 sg13g2_inv_1 _10369_ (.Y(_04375_),
    .A(_00088_));
 sg13g2_a21oi_1 _10370_ (.A1(net975),
    .A2(_04375_),
    .Y(_04376_),
    .B1(net1158));
 sg13g2_mux2_1 _10371_ (.A0(_00090_),
    .A1(_00091_),
    .S(net1221),
    .X(_04377_));
 sg13g2_a21o_1 _10372_ (.A2(_04377_),
    .A1(net1158),
    .B1(net1110),
    .X(_04378_));
 sg13g2_a21o_1 _10373_ (.A2(_04376_),
    .A1(_04374_),
    .B1(_04378_),
    .X(_04379_));
 sg13g2_mux4_1 _10374_ (.S0(net1158),
    .A0(_00092_),
    .A1(_00094_),
    .A2(_00093_),
    .A3(_00095_),
    .S1(net1221),
    .X(_04380_));
 sg13g2_inv_1 _10375_ (.Y(_04381_),
    .A(_04380_));
 sg13g2_a21oi_1 _10376_ (.A1(net1110),
    .A2(_04381_),
    .Y(_04382_),
    .B1(_03925_));
 sg13g2_inv_1 _10377_ (.Y(_04383_),
    .A(_00085_));
 sg13g2_o21ai_1 _10378_ (.B1(_04383_),
    .Y(_04384_),
    .A1(net1032),
    .A2(net1018));
 sg13g2_mux4_1 _10379_ (.S0(net1158),
    .A0(_00084_),
    .A1(_00086_),
    .A2(_04384_),
    .A3(_00087_),
    .S1(net1221),
    .X(_04385_));
 sg13g2_mux4_1 _10380_ (.S0(net1158),
    .A0(_00080_),
    .A1(_00082_),
    .A2(_00081_),
    .A3(_00083_),
    .S1(net1221),
    .X(_04386_));
 sg13g2_a21o_1 _10381_ (.A2(_04386_),
    .A1(net965),
    .B1(net946),
    .X(_04387_));
 sg13g2_a221oi_1 _10382_ (.B2(_04385_),
    .C1(_04387_),
    .B1(net968),
    .A1(_04379_),
    .Y(_04388_),
    .A2(_04382_));
 sg13g2_a21oi_2 _10383_ (.B1(_04388_),
    .Y(_04389_),
    .A2(_04372_),
    .A1(_04368_));
 sg13g2_buf_1 fanout744 (.A(net745),
    .X(net744));
 sg13g2_inv_2 _10385_ (.Y(_04391_),
    .A(net1253));
 sg13g2_o21ai_1 _10386_ (.B1(_04104_),
    .Y(_04392_),
    .A1(_04391_),
    .A2(net933));
 sg13g2_buf_2 fanout743 (.A(net745),
    .X(net743));
 sg13g2_nor2_1 _10388_ (.A(net906),
    .B(_04392_),
    .Y(_04394_));
 sg13g2_a21oi_1 _10389_ (.A1(_03389_),
    .A2(net906),
    .Y(_04395_),
    .B1(_04394_));
 sg13g2_xnor2_1 _10390_ (.Y(_04396_),
    .A(net872),
    .B(_04395_));
 sg13g2_buf_2 fanout742 (.A(net748),
    .X(net742));
 sg13g2_xnor2_1 _10392_ (.Y(_04398_),
    .A(_04389_),
    .B(_04396_));
 sg13g2_nand3_1 _10393_ (.B(_04353_),
    .C(_04398_),
    .A(_04350_),
    .Y(_04399_));
 sg13g2_nor2_1 _10394_ (.A(_04289_),
    .B(_04399_),
    .Y(_04400_));
 sg13g2_mux2_1 _10395_ (.A0(_00495_),
    .A1(_00497_),
    .S(net1161),
    .X(_04401_));
 sg13g2_a221oi_1 _10396_ (.B2(net1223),
    .C1(net1110),
    .B1(_04401_),
    .A1(_00496_),
    .Y(_04402_),
    .A2(_04238_));
 sg13g2_mux4_1 _10397_ (.S0(net1161),
    .A0(_00498_),
    .A1(_00500_),
    .A2(_00499_),
    .A3(_00501_),
    .S1(net1223),
    .X(_04403_));
 sg13g2_o21ai_1 _10398_ (.B1(net1002),
    .Y(_04404_),
    .A1(net961),
    .A2(_04403_));
 sg13g2_or2_1 _10399_ (.X(_04405_),
    .B(_04404_),
    .A(_04402_));
 sg13g2_mux4_1 _10400_ (.S0(net1160),
    .A0(_00502_),
    .A1(_00504_),
    .A2(_00503_),
    .A3(_00505_),
    .S1(net1222),
    .X(_04406_));
 sg13g2_and2_1 _10401_ (.A(net992),
    .B(_04406_),
    .X(_04407_));
 sg13g2_mux4_1 _10402_ (.S0(net1160),
    .A0(_00506_),
    .A1(_00508_),
    .A2(_00507_),
    .A3(_00509_),
    .S1(net1222),
    .X(_04408_));
 sg13g2_and2_1 _10403_ (.A(net969),
    .B(_04408_),
    .X(_04409_));
 sg13g2_or2_2 _10404_ (.X(_04410_),
    .B(net1107),
    .A(net1139));
 sg13g2_buf_2 fanout741 (.A(net742),
    .X(net741));
 sg13g2_o21ai_1 _10406_ (.B1(_00494_),
    .Y(_04412_),
    .A1(net975),
    .A2(_00495_));
 sg13g2_nor3_1 _10407_ (.A(net1398),
    .B(_04410_),
    .C(_04412_),
    .Y(_04413_));
 sg13g2_nor4_2 _10408_ (.A(net946),
    .B(_04407_),
    .C(_04409_),
    .Y(_04414_),
    .D(_04413_));
 sg13g2_mux4_1 _10409_ (.S0(net1160),
    .A0(_00486_),
    .A1(_00488_),
    .A2(_00487_),
    .A3(_00489_),
    .S1(net1222),
    .X(_04415_));
 sg13g2_and2_1 _10410_ (.A(net991),
    .B(_04415_),
    .X(_04416_));
 sg13g2_mux4_1 _10411_ (.S0(net1160),
    .A0(_00490_),
    .A1(_00492_),
    .A2(_00491_),
    .A3(_00493_),
    .S1(net1222),
    .X(_04417_));
 sg13g2_nand2_1 _10412_ (.Y(_04418_),
    .A(net1398),
    .B(_04417_));
 sg13g2_mux4_1 _10413_ (.S0(net1160),
    .A0(_00482_),
    .A1(_00484_),
    .A2(_00483_),
    .A3(_00485_),
    .S1(net1222),
    .X(_04419_));
 sg13g2_nand2_1 _10414_ (.Y(_04420_),
    .A(net1002),
    .B(_04419_));
 sg13g2_a21oi_1 _10415_ (.A1(_04418_),
    .A2(_04420_),
    .Y(_04421_),
    .B1(net961));
 sg13g2_nand2_1 _10416_ (.Y(_04422_),
    .A(net1143),
    .B(_00480_));
 sg13g2_nor2b_1 _10417_ (.A(net1143),
    .B_N(_00479_),
    .Y(_04423_));
 sg13g2_a22oi_1 _10418_ (.Y(_04424_),
    .B1(_04423_),
    .B2(net973),
    .A2(_00481_),
    .A1(net1143));
 sg13g2_a22oi_1 _10419_ (.Y(_04425_),
    .B1(_04424_),
    .B2(_04245_),
    .A2(_04422_),
    .A1(net972));
 sg13g2_nor4_2 _10420_ (.A(_04141_),
    .B(_04416_),
    .C(_04421_),
    .Y(_04426_),
    .D(_04425_));
 sg13g2_a21o_2 _10421_ (.A2(_04414_),
    .A1(_04405_),
    .B1(_04426_),
    .X(_04427_));
 sg13g2_buf_2 fanout740 (.A(net748),
    .X(net740));
 sg13g2_or4_1 _10423_ (.A(net918),
    .B(_03826_),
    .C(_03828_),
    .D(_03830_),
    .X(_04429_));
 sg13g2_buf_2 fanout739 (.A(net748),
    .X(net739));
 sg13g2_buf_1 fanout738 (.A(_08271_),
    .X(net738));
 sg13g2_nor4_1 _10426_ (.A(_03013_),
    .B(_03018_),
    .C(_03028_),
    .D(net903),
    .Y(_04432_));
 sg13g2_buf_2 fanout737 (.A(net738),
    .X(net737));
 sg13g2_nand4_1 _10428_ (.B(net1255),
    .C(_02561_),
    .A(net1252),
    .Y(_04434_),
    .D(_03824_));
 sg13g2_buf_2 fanout736 (.A(net738),
    .X(net736));
 sg13g2_nor2b_1 _10430_ (.A(_04104_),
    .B_N(_04434_),
    .Y(_04436_));
 sg13g2_buf_2 fanout735 (.A(net738),
    .X(net735));
 sg13g2_buf_1 fanout734 (.A(net735),
    .X(net734));
 sg13g2_a21oi_1 _10433_ (.A1(net933),
    .A2(_04434_),
    .Y(_04439_),
    .B1(net961));
 sg13g2_nor3_1 _10434_ (.A(net907),
    .B(net897),
    .C(_04439_),
    .Y(_04440_));
 sg13g2_a21oi_1 _10435_ (.A1(_03048_),
    .A2(_04432_),
    .Y(_04441_),
    .B1(_04440_));
 sg13g2_xnor2_1 _10436_ (.Y(_04442_),
    .A(net880),
    .B(_04441_));
 sg13g2_xnor2_1 _10437_ (.Y(_04443_),
    .A(_04427_),
    .B(_04442_));
 sg13g2_buf_2 fanout733 (.A(net735),
    .X(net733));
 sg13g2_nor2b_1 _10439_ (.A(_00473_),
    .B_N(net1163),
    .Y(_04445_));
 sg13g2_o21ai_1 _10440_ (.B1(_04445_),
    .Y(_04446_),
    .A1(net1035),
    .A2(net1021));
 sg13g2_o21ai_1 _10441_ (.B1(_04446_),
    .Y(_04447_),
    .A1(net1163),
    .A2(_00471_));
 sg13g2_buf_1 fanout732 (.A(_08271_),
    .X(net732));
 sg13g2_buf_2 fanout731 (.A(net732),
    .X(net731));
 sg13g2_nor2b_1 _10444_ (.A(net1163),
    .B_N(_00476_),
    .Y(_04450_));
 sg13g2_a22oi_1 _10445_ (.Y(_04451_),
    .B1(net1006),
    .B2(_04450_),
    .A2(_00478_),
    .A1(net1163));
 sg13g2_nor2b_1 _10446_ (.A(net1163),
    .B_N(_00475_),
    .Y(_04452_));
 sg13g2_a22oi_1 _10447_ (.Y(_04453_),
    .B1(net1007),
    .B2(_04452_),
    .A2(_00477_),
    .A1(net1163));
 sg13g2_nor2b_1 _10448_ (.A(net1163),
    .B_N(_00472_),
    .Y(_04454_));
 sg13g2_a22oi_1 _10449_ (.Y(_04455_),
    .B1(net1004),
    .B2(_04454_),
    .A2(_00474_),
    .A1(net1163));
 sg13g2_or3_1 _10450_ (.A(_04451_),
    .B(_04453_),
    .C(_04455_),
    .X(_04456_));
 sg13g2_o21ai_1 _10451_ (.B1(net993),
    .Y(_04457_),
    .A1(net1038),
    .A2(net1023));
 sg13g2_buf_2 fanout730 (.A(net732),
    .X(net730));
 sg13g2_buf_1 fanout729 (.A(net730),
    .X(net729));
 sg13g2_a22oi_1 _10454_ (.Y(_04460_),
    .B1(_04456_),
    .B2(net916),
    .A2(_04447_),
    .A1(net1040));
 sg13g2_nor2b_1 _10455_ (.A(net1165),
    .B_N(_00456_),
    .Y(_04461_));
 sg13g2_a22oi_1 _10456_ (.Y(_04462_),
    .B1(net1004),
    .B2(_04461_),
    .A2(_00458_),
    .A1(net1165));
 sg13g2_mux4_1 _10457_ (.S0(net1164),
    .A0(_00459_),
    .A1(_00461_),
    .A2(_00460_),
    .A3(_00462_),
    .S1(net1225),
    .X(_04463_));
 sg13g2_nor2_1 _10458_ (.A(net962),
    .B(_04463_),
    .Y(_04464_));
 sg13g2_or3_1 _10459_ (.A(net947),
    .B(_04462_),
    .C(_04464_),
    .X(_04465_));
 sg13g2_or2_1 _10460_ (.X(_04466_),
    .B(_00455_),
    .A(net1140));
 sg13g2_nor2b_1 _10461_ (.A(_00457_),
    .B_N(net1165),
    .Y(_04467_));
 sg13g2_o21ai_1 _10462_ (.B1(_04467_),
    .Y(_04468_),
    .A1(net1035),
    .A2(net1021));
 sg13g2_a21oi_1 _10463_ (.A1(_04466_),
    .A2(_04468_),
    .Y(_04469_),
    .B1(net998));
 sg13g2_mux4_1 _10464_ (.S0(net1138),
    .A0(_00467_),
    .A1(_00469_),
    .A2(_00468_),
    .A3(_00470_),
    .S1(net1212),
    .X(_04470_));
 sg13g2_mux4_1 _10465_ (.S0(net1138),
    .A0(_00451_),
    .A1(_00453_),
    .A2(_00452_),
    .A3(_00454_),
    .S1(net1212),
    .X(_04471_));
 sg13g2_nor2_1 _10466_ (.A(net1393),
    .B(_03735_),
    .Y(_04472_));
 sg13g2_a221oi_1 _10467_ (.B2(_04472_),
    .C1(net920),
    .B1(_04471_),
    .A1(net925),
    .Y(_04473_),
    .A2(_04470_));
 sg13g2_o21ai_1 _10468_ (.B1(_04473_),
    .Y(_04474_),
    .A1(_04465_),
    .A2(_04469_));
 sg13g2_nor2b_1 _10469_ (.A(net1165),
    .B_N(_00448_),
    .Y(_04475_));
 sg13g2_a22oi_1 _10470_ (.Y(_04476_),
    .B1(_04475_),
    .B2(net976),
    .A2(_00450_),
    .A1(net1165));
 sg13g2_nand2b_2 _10471_ (.Y(_04477_),
    .B(net1144),
    .A_N(net1214));
 sg13g2_buf_2 fanout728 (.A(net730),
    .X(net728));
 sg13g2_buf_2 fanout727 (.A(_08350_),
    .X(net727));
 sg13g2_o21ai_1 _10474_ (.B1(net994),
    .Y(_04480_),
    .A1(_00449_),
    .A2(_04477_));
 sg13g2_nor2_1 _10475_ (.A(net995),
    .B(_04245_),
    .Y(_04481_));
 sg13g2_buf_2 fanout726 (.A(net727),
    .X(net726));
 sg13g2_mux4_1 _10477_ (.S0(net1165),
    .A0(_00463_),
    .A1(_00465_),
    .A2(_00464_),
    .A3(_00466_),
    .S1(net1225),
    .X(_04483_));
 sg13g2_nand3_1 _10478_ (.B(net915),
    .C(_04483_),
    .A(net935),
    .Y(_04484_));
 sg13g2_o21ai_1 _10479_ (.B1(_04484_),
    .Y(_04485_),
    .A1(_04476_),
    .A2(_04480_));
 sg13g2_or3_1 _10480_ (.A(_04460_),
    .B(_04474_),
    .C(_04485_),
    .X(_04486_));
 sg13g2_buf_2 fanout725 (.A(net727),
    .X(net725));
 sg13g2_nand2_2 _10482_ (.Y(_04488_),
    .A(net940),
    .B(_04434_));
 sg13g2_buf_2 fanout724 (.A(net727),
    .X(net724));
 sg13g2_a21oi_2 _10484_ (.B1(net897),
    .Y(_04490_),
    .A2(net896),
    .A1(net1398));
 sg13g2_nor2_1 _10485_ (.A(net907),
    .B(_04490_),
    .Y(_04491_));
 sg13g2_nor3_1 _10486_ (.A(net949),
    .B(_03078_),
    .C(net900),
    .Y(_04492_));
 sg13g2_nor3_1 _10487_ (.A(net880),
    .B(_04491_),
    .C(_04492_),
    .Y(_04493_));
 sg13g2_nand2b_1 _10488_ (.Y(_04494_),
    .B(net900),
    .A_N(_04490_));
 sg13g2_or3_1 _10489_ (.A(net950),
    .B(_03078_),
    .C(net899),
    .X(_04495_));
 sg13g2_a21oi_1 _10490_ (.A1(_04494_),
    .A2(_04495_),
    .Y(_04496_),
    .B1(net873));
 sg13g2_nor3_2 _10491_ (.A(net625),
    .B(_04493_),
    .C(_04496_),
    .Y(_04497_));
 sg13g2_buf_2 fanout723 (.A(net727),
    .X(net723));
 sg13g2_buf_1 fanout722 (.A(_08350_),
    .X(net722));
 sg13g2_nand3_1 _10494_ (.B(_04494_),
    .C(_04495_),
    .A(net873),
    .Y(_04500_));
 sg13g2_o21ai_1 _10495_ (.B1(net880),
    .Y(_04501_),
    .A1(_04491_),
    .A2(_04492_));
 sg13g2_inv_1 _10496_ (.Y(_04502_),
    .A(net624));
 sg13g2_a21oi_2 _10497_ (.B1(_04502_),
    .Y(_04503_),
    .A2(_04501_),
    .A1(_04500_));
 sg13g2_nor2_1 _10498_ (.A(_04497_),
    .B(_04503_),
    .Y(_04504_));
 sg13g2_a21oi_2 _10499_ (.B1(net897),
    .Y(_04505_),
    .A2(net896),
    .A1(net1162));
 sg13g2_mux2_1 _10500_ (.A0(_03007_),
    .A1(_04505_),
    .S(net900),
    .X(_04506_));
 sg13g2_xnor2_1 _10501_ (.Y(_04507_),
    .A(net873),
    .B(_04506_));
 sg13g2_nor2_1 _10502_ (.A(net959),
    .B(_00536_),
    .Y(_04508_));
 sg13g2_nor2_1 _10503_ (.A(net1168),
    .B(_00534_),
    .Y(_04509_));
 sg13g2_a21oi_1 _10504_ (.A1(net935),
    .A2(_04508_),
    .Y(_04510_),
    .B1(_04509_));
 sg13g2_mux4_1 _10505_ (.S0(net1168),
    .A0(_00535_),
    .A1(_00537_),
    .A2(_00539_),
    .A3(_00541_),
    .S1(net1113),
    .X(_04511_));
 sg13g2_inv_1 _10506_ (.Y(_04512_),
    .A(_04511_));
 sg13g2_buf_2 fanout721 (.A(net722),
    .X(net721));
 sg13g2_nor2b_1 _10508_ (.A(net1167),
    .B_N(_00538_),
    .Y(_04514_));
 sg13g2_a22oi_1 _10509_ (.Y(_04515_),
    .B1(net1008),
    .B2(_04514_),
    .A2(_00540_),
    .A1(net1169));
 sg13g2_a22oi_1 _10510_ (.Y(_04516_),
    .B1(_04515_),
    .B2(net916),
    .A2(_04512_),
    .A1(net1225));
 sg13g2_o21ai_1 _10511_ (.B1(_04516_),
    .Y(_04517_),
    .A1(net998),
    .A2(_04510_));
 sg13g2_o21ai_1 _10512_ (.B1(_03935_),
    .Y(_04518_),
    .A1(net1034),
    .A2(net1023));
 sg13g2_buf_2 fanout720 (.A(net721),
    .X(net720));
 sg13g2_nor2b_1 _10514_ (.A(net1182),
    .B_N(_00522_),
    .Y(_04520_));
 sg13g2_a22oi_1 _10515_ (.Y(_04521_),
    .B1(_04518_),
    .B2(_04520_),
    .A2(_00524_),
    .A1(net1182));
 sg13g2_mux4_1 _10516_ (.S0(net1182),
    .A0(_00519_),
    .A1(_00521_),
    .A2(_00523_),
    .A3(_00525_),
    .S1(net1113),
    .X(_04522_));
 sg13g2_nor2_1 _10517_ (.A(net976),
    .B(_04522_),
    .Y(_04523_));
 sg13g2_or2_1 _10518_ (.X(_04524_),
    .B(_00518_),
    .A(net1175));
 sg13g2_nor2b_1 _10519_ (.A(_00520_),
    .B_N(net1175),
    .Y(_04525_));
 sg13g2_o21ai_1 _10520_ (.B1(_04525_),
    .Y(_04526_),
    .A1(net1035),
    .A2(net1021));
 sg13g2_a21oi_1 _10521_ (.A1(_04524_),
    .A2(_04526_),
    .Y(_04527_),
    .B1(net999));
 sg13g2_or4_1 _10522_ (.A(net947),
    .B(_04521_),
    .C(_04523_),
    .D(_04527_),
    .X(_04528_));
 sg13g2_buf_2 fanout719 (.A(net722),
    .X(net719));
 sg13g2_nand2_1 _10524_ (.Y(_04530_),
    .A(_00511_),
    .B(_00510_));
 sg13g2_a22oi_1 _10525_ (.Y(_04531_),
    .B1(_04410_),
    .B2(net988),
    .A2(_04530_),
    .A1(net1227));
 sg13g2_nand2_1 _10526_ (.Y(_04532_),
    .A(net1178),
    .B(_00517_));
 sg13g2_nand2b_1 _10527_ (.Y(_04533_),
    .B(_00515_),
    .A_N(net1178));
 sg13g2_a22oi_1 _10528_ (.Y(_04534_),
    .B1(net1006),
    .B2(net988),
    .A2(_04533_),
    .A1(_04532_));
 sg13g2_nand2_1 _10529_ (.Y(_04535_),
    .A(net1178),
    .B(_00516_));
 sg13g2_nand2b_1 _10530_ (.Y(_04536_),
    .B(_00514_),
    .A_N(net1178));
 sg13g2_a22oi_1 _10531_ (.Y(_04537_),
    .B1(net1008),
    .B2(net988),
    .A2(_04536_),
    .A1(_04535_));
 sg13g2_nor4_1 _10532_ (.A(net921),
    .B(_04531_),
    .C(_04534_),
    .D(_04537_),
    .Y(_04538_));
 sg13g2_mux4_1 _10533_ (.S0(net1169),
    .A0(_00530_),
    .A1(_00532_),
    .A2(_00531_),
    .A3(_00533_),
    .S1(net1225),
    .X(_04539_));
 sg13g2_nand2_1 _10534_ (.Y(_04540_),
    .A(net925),
    .B(_04539_));
 sg13g2_nand2_1 _10535_ (.Y(_04541_),
    .A(net1169),
    .B(_00513_));
 sg13g2_nand2b_1 _10536_ (.Y(_04542_),
    .B(_00511_),
    .A_N(net1169));
 sg13g2_a21oi_1 _10537_ (.A1(_04541_),
    .A2(_04542_),
    .Y(_04543_),
    .B1(net976));
 sg13g2_and2_1 _10538_ (.A(_00512_),
    .B(_04238_),
    .X(_04544_));
 sg13g2_o21ai_1 _10539_ (.B1(net994),
    .Y(_04545_),
    .A1(_04543_),
    .A2(_04544_));
 sg13g2_mux4_1 _10540_ (.S0(net1168),
    .A0(_00526_),
    .A1(_00528_),
    .A2(_00527_),
    .A3(_00529_),
    .S1(net1225),
    .X(_04546_));
 sg13g2_nand2_1 _10541_ (.Y(_04547_),
    .A(net914),
    .B(_04546_));
 sg13g2_and4_1 _10542_ (.A(_04538_),
    .B(_04540_),
    .C(_04545_),
    .D(_04547_),
    .X(_04548_));
 sg13g2_buf_2 fanout718 (.A(net722),
    .X(net718));
 sg13g2_nand3_1 _10544_ (.B(_04528_),
    .C(_04548_),
    .A(_04517_),
    .Y(_04550_));
 sg13g2_buf_2 fanout717 (.A(_08429_),
    .X(net717));
 sg13g2_nor2_1 _10546_ (.A(_04507_),
    .B(_04550_),
    .Y(_04552_));
 sg13g2_and2_1 _10547_ (.A(_04507_),
    .B(_04550_),
    .X(_04553_));
 sg13g2_nor2_1 _10548_ (.A(_04552_),
    .B(_04553_),
    .Y(_04554_));
 sg13g2_nor2b_1 _10549_ (.A(_00425_),
    .B_N(net1140),
    .Y(_04555_));
 sg13g2_o21ai_1 _10550_ (.B1(_04555_),
    .Y(_04556_),
    .A1(net1028),
    .A2(net1014));
 sg13g2_o21ai_1 _10551_ (.B1(_04556_),
    .Y(_04557_),
    .A1(net1140),
    .A2(_00423_));
 sg13g2_nor2b_1 _10552_ (.A(net1139),
    .B_N(_00424_),
    .Y(_04558_));
 sg13g2_a22oi_1 _10553_ (.Y(_04559_),
    .B1(net1004),
    .B2(_04558_),
    .A2(_00426_),
    .A1(net1139));
 sg13g2_mux4_1 _10554_ (.S0(net1138),
    .A0(_00427_),
    .A1(_00429_),
    .A2(_00428_),
    .A3(_00430_),
    .S1(net1212),
    .X(_04560_));
 sg13g2_nor2_1 _10555_ (.A(net961),
    .B(_04560_),
    .Y(_04561_));
 sg13g2_or2_1 _10556_ (.X(_04562_),
    .B(_04561_),
    .A(_04559_));
 sg13g2_a22oi_1 _10557_ (.Y(_04563_),
    .B1(_04562_),
    .B2(net947),
    .A2(_04557_),
    .A1(net1040));
 sg13g2_mux4_1 _10558_ (.S0(net1144),
    .A0(_00435_),
    .A1(_00437_),
    .A2(_00436_),
    .A3(_00438_),
    .S1(net1214),
    .X(_04564_));
 sg13g2_nand2_1 _10559_ (.Y(_04565_),
    .A(net1392),
    .B(_04564_));
 sg13g2_mux2_1 _10560_ (.A0(_00420_),
    .A1(_00422_),
    .S(net1145),
    .X(_04566_));
 sg13g2_nand3_1 _10561_ (.B(net995),
    .C(_04566_),
    .A(net1214),
    .Y(_04567_));
 sg13g2_a21oi_1 _10562_ (.A1(_04565_),
    .A2(_04567_),
    .Y(_04568_),
    .B1(_03735_));
 sg13g2_o21ai_1 _10563_ (.B1(net994),
    .Y(_04569_),
    .A1(_00417_),
    .A2(_04477_));
 sg13g2_mux2_1 _10564_ (.A0(_00431_),
    .A1(_00433_),
    .S(net1140),
    .X(_04570_));
 sg13g2_nand3_1 _10565_ (.B(net965),
    .C(_04570_),
    .A(net1393),
    .Y(_04571_));
 sg13g2_mux2_1 _10566_ (.A0(_00416_),
    .A1(_00418_),
    .S(net1145),
    .X(_04572_));
 sg13g2_a21oi_1 _10567_ (.A1(net994),
    .A2(_04572_),
    .Y(_04573_),
    .B1(net972));
 sg13g2_a21oi_1 _10568_ (.A1(_04569_),
    .A2(_04571_),
    .Y(_04574_),
    .B1(_04573_));
 sg13g2_mux2_1 _10569_ (.A0(_00432_),
    .A1(_00434_),
    .S(net1145),
    .X(_04575_));
 sg13g2_nand4_1 _10570_ (.B(net1393),
    .C(net965),
    .A(net1214),
    .Y(_04576_),
    .D(_04575_));
 sg13g2_nor2_2 _10571_ (.A(net1399),
    .B(net1394),
    .Y(_04577_));
 sg13g2_buf_2 fanout716 (.A(net717),
    .X(net716));
 sg13g2_mux2_1 _10573_ (.A0(_00419_),
    .A1(_00421_),
    .S(net1145),
    .X(_04579_));
 sg13g2_nand3_1 _10574_ (.B(_04577_),
    .C(_04579_),
    .A(_03935_),
    .Y(_04580_));
 sg13g2_nand3_1 _10575_ (.B(_04576_),
    .C(_04580_),
    .A(net928),
    .Y(_04581_));
 sg13g2_or3_1 _10576_ (.A(_04568_),
    .B(_04574_),
    .C(_04581_),
    .X(_04582_));
 sg13g2_mux4_1 _10577_ (.S0(net1139),
    .A0(_00440_),
    .A1(_00442_),
    .A2(_00444_),
    .A3(_00446_),
    .S1(net1107),
    .X(_04583_));
 sg13g2_nor2_1 _10578_ (.A(net972),
    .B(_04583_),
    .Y(_04584_));
 sg13g2_nor2b_1 _10579_ (.A(net1139),
    .B_N(_00443_),
    .Y(_04585_));
 sg13g2_a22oi_1 _10580_ (.Y(_04586_),
    .B1(net1007),
    .B2(_04585_),
    .A2(_00445_),
    .A1(net1140));
 sg13g2_inv_1 _10581_ (.Y(_04587_),
    .A(_00441_));
 sg13g2_o21ai_1 _10582_ (.B1(_04587_),
    .Y(_04588_),
    .A1(net1029),
    .A2(net1015));
 sg13g2_nor2b_1 _10583_ (.A(net1140),
    .B_N(_00439_),
    .Y(_04589_));
 sg13g2_a22oi_1 _10584_ (.Y(_04590_),
    .B1(_04589_),
    .B2(net1001),
    .A2(_04588_),
    .A1(net1140));
 sg13g2_nor4_1 _10585_ (.A(net916),
    .B(_04584_),
    .C(_04586_),
    .D(_04590_),
    .Y(_04591_));
 sg13g2_or3_1 _10586_ (.A(_04563_),
    .B(_04582_),
    .C(_04591_),
    .X(_04592_));
 sg13g2_buf_2 fanout715 (.A(net716),
    .X(net715));
 sg13g2_and2_1 _10588_ (.A(_03080_),
    .B(net907),
    .X(_04594_));
 sg13g2_a22oi_1 _10589_ (.Y(_04595_),
    .B1(net897),
    .B2(net907),
    .A2(net896),
    .A1(net1395));
 sg13g2_a21oi_1 _10590_ (.A1(_03109_),
    .A2(_04594_),
    .Y(_04596_),
    .B1(_04595_));
 sg13g2_xnor2_1 _10591_ (.Y(_04597_),
    .A(net873),
    .B(_04596_));
 sg13g2_xnor2_1 _10592_ (.Y(_04598_),
    .A(_04592_),
    .B(_04597_));
 sg13g2_buf_2 fanout714 (.A(net717),
    .X(net714));
 sg13g2_nand4_1 _10594_ (.B(_04504_),
    .C(_04554_),
    .A(_04443_),
    .Y(_04600_),
    .D(_04598_));
 sg13g2_buf_2 fanout713 (.A(net717),
    .X(net713));
 sg13g2_or2_1 _10596_ (.X(_04602_),
    .B(_00336_),
    .A(net1155));
 sg13g2_nor2b_1 _10597_ (.A(_00338_),
    .B_N(net1158),
    .Y(_04603_));
 sg13g2_o21ai_1 _10598_ (.B1(_04603_),
    .Y(_04604_),
    .A1(net1031),
    .A2(net1017));
 sg13g2_a21oi_1 _10599_ (.A1(_04602_),
    .A2(_04604_),
    .Y(_04605_),
    .B1(net1217));
 sg13g2_mux2_1 _10600_ (.A0(_00337_),
    .A1(_00339_),
    .S(net1155),
    .X(_04606_));
 sg13g2_o21ai_1 _10601_ (.B1(net965),
    .Y(_04607_),
    .A1(net974),
    .A2(_04606_));
 sg13g2_nor3_1 _10602_ (.A(_00336_),
    .B(net1031),
    .C(net1017),
    .Y(_04608_));
 sg13g2_a21o_1 _10603_ (.A2(_04607_),
    .A1(net932),
    .B1(_04608_),
    .X(_04609_));
 sg13g2_mux4_1 _10604_ (.S0(net1155),
    .A0(_00340_),
    .A1(_00342_),
    .A2(_00341_),
    .A3(_00343_),
    .S1(net1217),
    .X(_04610_));
 sg13g2_and2_1 _10605_ (.A(net968),
    .B(_04610_),
    .X(_04611_));
 sg13g2_mux4_1 _10606_ (.S0(net1155),
    .A0(_00348_),
    .A1(_00350_),
    .A2(_00349_),
    .A3(_00351_),
    .S1(net1218),
    .X(_04612_));
 sg13g2_and2_1 _10607_ (.A(net969),
    .B(_04612_),
    .X(_04613_));
 sg13g2_mux4_1 _10608_ (.S0(net1155),
    .A0(_00344_),
    .A1(_00346_),
    .A2(_00345_),
    .A3(_00347_),
    .S1(net1218),
    .X(_04614_));
 sg13g2_and2_1 _10609_ (.A(net991),
    .B(_04614_),
    .X(_04615_));
 sg13g2_nor4_1 _10610_ (.A(net946),
    .B(_04611_),
    .C(_04613_),
    .D(_04615_),
    .Y(_04616_));
 sg13g2_o21ai_1 _10611_ (.B1(_04616_),
    .Y(_04617_),
    .A1(_04605_),
    .A2(_04609_));
 sg13g2_or2_1 _10612_ (.X(_04618_),
    .B(_00320_),
    .A(net1156));
 sg13g2_nor2b_1 _10613_ (.A(_00322_),
    .B_N(net1156),
    .Y(_04619_));
 sg13g2_o21ai_1 _10614_ (.B1(_04619_),
    .Y(_04620_),
    .A1(net1032),
    .A2(net1018));
 sg13g2_a21oi_1 _10615_ (.A1(_04618_),
    .A2(_04620_),
    .Y(_04621_),
    .B1(net1220));
 sg13g2_mux2_1 _10616_ (.A0(_00321_),
    .A1(_00323_),
    .S(net1157),
    .X(_04622_));
 sg13g2_o21ai_1 _10617_ (.B1(net964),
    .Y(_04623_),
    .A1(net974),
    .A2(_04622_));
 sg13g2_nor3_1 _10618_ (.A(_00320_),
    .B(net1030),
    .C(net1016),
    .Y(_04624_));
 sg13g2_a21o_1 _10619_ (.A2(_04623_),
    .A1(net932),
    .B1(_04624_),
    .X(_04625_));
 sg13g2_mux4_1 _10620_ (.S0(net1156),
    .A0(_00328_),
    .A1(_00330_),
    .A2(_00329_),
    .A3(_00331_),
    .S1(net1219),
    .X(_04626_));
 sg13g2_mux4_1 _10621_ (.S0(net1150),
    .A0(_00324_),
    .A1(_00326_),
    .A2(_00325_),
    .A3(_00327_),
    .S1(net1219),
    .X(_04627_));
 sg13g2_mux4_1 _10622_ (.S0(net1150),
    .A0(_00332_),
    .A1(_00334_),
    .A2(_00333_),
    .A3(_00335_),
    .S1(net1219),
    .X(_04628_));
 sg13g2_mux4_1 _10623_ (.S0(net1398),
    .A0(_03743_),
    .A1(_04626_),
    .A2(_04627_),
    .A3(_04628_),
    .S1(net1110),
    .X(_04629_));
 sg13g2_nor2_1 _10624_ (.A(_03951_),
    .B(_04629_),
    .Y(_04630_));
 sg13g2_o21ai_1 _10625_ (.B1(_04630_),
    .Y(_04631_),
    .A1(_04621_),
    .A2(_04625_));
 sg13g2_nand2_1 _10626_ (.Y(_04632_),
    .A(_04617_),
    .B(_04631_));
 sg13g2_buf_2 fanout712 (.A(net717),
    .X(net712));
 sg13g2_a22oi_1 _10628_ (.Y(_04634_),
    .B1(net900),
    .B2(_03817_),
    .A2(_03810_),
    .A1(_03805_));
 sg13g2_o21ai_1 _10629_ (.B1(_04634_),
    .Y(_04635_),
    .A1(net949),
    .A2(_03206_));
 sg13g2_a21oi_2 _10630_ (.B1(_03893_),
    .Y(_04636_),
    .A2(net918),
    .A1(net1276));
 sg13g2_or3_1 _10631_ (.A(net878),
    .B(net904),
    .C(_04636_),
    .X(_04637_));
 sg13g2_nand3_1 _10632_ (.B(net899),
    .C(_04636_),
    .A(net878),
    .Y(_04638_));
 sg13g2_or4_1 _10633_ (.A(net949),
    .B(_03206_),
    .C(net878),
    .D(net899),
    .X(_04639_));
 sg13g2_nand4_1 _10634_ (.B(_04637_),
    .C(_04638_),
    .A(_04635_),
    .Y(_04640_),
    .D(_04639_));
 sg13g2_buf_2 fanout711 (.A(net712),
    .X(net711));
 sg13g2_xnor2_1 _10636_ (.Y(_04642_),
    .A(net621),
    .B(_04640_));
 sg13g2_or2_1 _10637_ (.X(_04643_),
    .B(_00304_),
    .A(net1211));
 sg13g2_nor2b_1 _10638_ (.A(_00305_),
    .B_N(net1211),
    .Y(_04644_));
 sg13g2_o21ai_1 _10639_ (.B1(_04644_),
    .Y(_04645_),
    .A1(net1028),
    .A2(net1014));
 sg13g2_a21o_1 _10640_ (.A2(_04645_),
    .A1(_04643_),
    .B1(net1136),
    .X(_04646_));
 sg13g2_and2_1 _10641_ (.A(net1211),
    .B(_00307_),
    .X(_04647_));
 sg13g2_a22oi_1 _10642_ (.Y(_04648_),
    .B1(_04647_),
    .B2(net958),
    .A2(_00306_),
    .A1(net970));
 sg13g2_o21ai_1 _10643_ (.B1(net926),
    .Y(_04649_),
    .A1(_04245_),
    .A2(_04648_));
 sg13g2_nand2b_1 _10644_ (.Y(_04650_),
    .B(net920),
    .A_N(_00304_));
 sg13g2_nand3_1 _10645_ (.B(_04649_),
    .C(_04650_),
    .A(_04646_),
    .Y(_04651_));
 sg13g2_mux4_1 _10646_ (.S0(net1135),
    .A0(_00316_),
    .A1(_00318_),
    .A2(_00317_),
    .A3(_00319_),
    .S1(net1211),
    .X(_04652_));
 sg13g2_mux2_1 _10647_ (.A0(_00313_),
    .A1(_00315_),
    .S(net1136),
    .X(_04653_));
 sg13g2_nand2b_1 _10648_ (.Y(_04654_),
    .B(_04653_),
    .A_N(_04045_));
 sg13g2_mux2_1 _10649_ (.A0(_00309_),
    .A1(_00311_),
    .S(net1135),
    .X(_04655_));
 sg13g2_nand3_1 _10650_ (.B(net967),
    .C(_04655_),
    .A(net1211),
    .Y(_04656_));
 sg13g2_mux2_1 _10651_ (.A0(_00312_),
    .A1(_00314_),
    .S(net1135),
    .X(_04657_));
 sg13g2_nand3_1 _10652_ (.B(net1040),
    .C(_04657_),
    .A(net1397),
    .Y(_04658_));
 sg13g2_mux2_1 _10653_ (.A0(_00308_),
    .A1(_00310_),
    .S(net1135),
    .X(_04659_));
 sg13g2_nand3_1 _10654_ (.B(net967),
    .C(_04659_),
    .A(net970),
    .Y(_04660_));
 sg13g2_nand4_1 _10655_ (.B(_04656_),
    .C(_04658_),
    .A(_04654_),
    .Y(_04661_),
    .D(_04660_));
 sg13g2_a22oi_1 _10656_ (.Y(_04662_),
    .B1(_04661_),
    .B2(net945),
    .A2(_04652_),
    .A1(_04144_));
 sg13g2_nor2b_1 _10657_ (.A(net1141),
    .B_N(_00300_),
    .Y(_04663_));
 sg13g2_a22oi_1 _10658_ (.Y(_04664_),
    .B1(net1007),
    .B2(_04663_),
    .A2(_00302_),
    .A1(net1141));
 sg13g2_nor2_1 _10659_ (.A(_00296_),
    .B(_03781_),
    .Y(_04665_));
 sg13g2_nor2_1 _10660_ (.A(_04664_),
    .B(_04665_),
    .Y(_04666_));
 sg13g2_nor2b_1 _10661_ (.A(net1108),
    .B_N(_00297_),
    .Y(_04667_));
 sg13g2_a22oi_1 _10662_ (.Y(_04668_),
    .B1(net990),
    .B2(_04667_),
    .A2(_00301_),
    .A1(net1108));
 sg13g2_nor3_1 _10663_ (.A(net1107),
    .B(_00298_),
    .C(_04477_),
    .Y(_04669_));
 sg13g2_nor2b_1 _10664_ (.A(net1107),
    .B_N(_00299_),
    .Y(_04670_));
 sg13g2_a22oi_1 _10665_ (.Y(_04671_),
    .B1(net987),
    .B2(_04670_),
    .A2(_00303_),
    .A1(net1107));
 sg13g2_nor4_1 _10666_ (.A(_03925_),
    .B(_04668_),
    .C(_04669_),
    .D(_04671_),
    .Y(_04672_));
 sg13g2_or2_1 _10667_ (.X(_04673_),
    .B(_00288_),
    .A(net1142));
 sg13g2_nor2b_1 _10668_ (.A(_00290_),
    .B_N(net1142),
    .Y(_04674_));
 sg13g2_o21ai_1 _10669_ (.B1(_04674_),
    .Y(_04675_),
    .A1(net1028),
    .A2(net1014));
 sg13g2_a21o_1 _10670_ (.A2(_04675_),
    .A1(_04673_),
    .B1(net1213),
    .X(_04676_));
 sg13g2_mux2_1 _10671_ (.A0(_00289_),
    .A1(_00291_),
    .S(net1142),
    .X(_04677_));
 sg13g2_o21ai_1 _10672_ (.B1(net963),
    .Y(_04678_),
    .A1(net972),
    .A2(_04677_));
 sg13g2_nor3_1 _10673_ (.A(_00288_),
    .B(net1028),
    .C(net1014),
    .Y(_04679_));
 sg13g2_a21oi_1 _10674_ (.A1(net928),
    .A2(_04678_),
    .Y(_04680_),
    .B1(_04679_));
 sg13g2_mux4_1 _10675_ (.S0(net1141),
    .A0(_00292_),
    .A1(_00294_),
    .A2(_00293_),
    .A3(_00295_),
    .S1(net1211),
    .X(_04681_));
 sg13g2_nand2_1 _10676_ (.Y(_04682_),
    .A(net967),
    .B(_04681_));
 sg13g2_nand3_1 _10677_ (.B(_04009_),
    .C(_04682_),
    .A(net928),
    .Y(_04683_));
 sg13g2_a221oi_1 _10678_ (.B2(_04680_),
    .C1(_04683_),
    .B1(_04676_),
    .A1(_04666_),
    .Y(_04684_),
    .A2(_04672_));
 sg13g2_a21o_2 _10679_ (.A2(_04662_),
    .A1(_04651_),
    .B1(_04684_),
    .X(_04685_));
 sg13g2_buf_2 fanout710 (.A(net711),
    .X(net710));
 sg13g2_a21oi_2 _10681_ (.B1(_03893_),
    .Y(_04687_),
    .A2(net918),
    .A1(net1265));
 sg13g2_mux2_1 _10682_ (.A0(_03236_),
    .A1(_04687_),
    .S(net899),
    .X(_04688_));
 sg13g2_xnor2_1 _10683_ (.Y(_04689_),
    .A(net878),
    .B(_04688_));
 sg13g2_xnor2_1 _10684_ (.Y(_04690_),
    .A(_04685_),
    .B(_04689_));
 sg13g2_mux4_1 _10685_ (.S0(net1129),
    .A0(_00364_),
    .A1(_00366_),
    .A2(_00365_),
    .A3(_00367_),
    .S1(net1207),
    .X(_04691_));
 sg13g2_mux4_1 _10686_ (.S0(net1130),
    .A0(_00360_),
    .A1(_00362_),
    .A2(_00361_),
    .A3(_00363_),
    .S1(net1207),
    .X(_04692_));
 sg13g2_mux2_1 _10687_ (.A0(_04691_),
    .A1(_04692_),
    .S(net961),
    .X(_04693_));
 sg13g2_mux4_1 _10688_ (.S0(net1129),
    .A0(_00356_),
    .A1(_00358_),
    .A2(_00357_),
    .A3(_00359_),
    .S1(net1207),
    .X(_04694_));
 sg13g2_and4_1 _10689_ (.A(net1109),
    .B(net1002),
    .C(net927),
    .D(_04694_),
    .X(_04695_));
 sg13g2_a22oi_1 _10690_ (.Y(_04696_),
    .B1(_04695_),
    .B2(_04141_),
    .A2(_04693_),
    .A1(net1397));
 sg13g2_or2_1 _10691_ (.X(_04697_),
    .B(_00352_),
    .A(net1131));
 sg13g2_nor2b_1 _10692_ (.A(_00354_),
    .B_N(net1131),
    .Y(_04698_));
 sg13g2_o21ai_1 _10693_ (.B1(_04698_),
    .Y(_04699_),
    .A1(net1027),
    .A2(net1013));
 sg13g2_a21o_1 _10694_ (.A2(_04699_),
    .A1(_04697_),
    .B1(net1209),
    .X(_04700_));
 sg13g2_nor2b_1 _10695_ (.A(net1128),
    .B_N(_00353_),
    .Y(_04701_));
 sg13g2_a22oi_1 _10696_ (.Y(_04702_),
    .B1(_04701_),
    .B2(net971),
    .A2(_00355_),
    .A1(net1128));
 sg13g2_o21ai_1 _10697_ (.B1(net927),
    .Y(_04703_),
    .A1(_04245_),
    .A2(_04702_));
 sg13g2_nand2b_1 _10698_ (.Y(_04704_),
    .B(net920),
    .A_N(_00352_));
 sg13g2_nand3_1 _10699_ (.B(_04703_),
    .C(_04704_),
    .A(_04700_),
    .Y(_04705_));
 sg13g2_or2_1 _10700_ (.X(_04706_),
    .B(_00368_),
    .A(net1128));
 sg13g2_nor2b_1 _10701_ (.A(_00370_),
    .B_N(net1128),
    .Y(_04707_));
 sg13g2_o21ai_1 _10702_ (.B1(_04707_),
    .Y(_04708_),
    .A1(net1025),
    .A2(net1011));
 sg13g2_a21o_1 _10703_ (.A2(_04708_),
    .A1(_04706_),
    .B1(net1207),
    .X(_04709_));
 sg13g2_mux2_1 _10704_ (.A0(_00369_),
    .A1(_00371_),
    .S(net1129),
    .X(_04710_));
 sg13g2_o21ai_1 _10705_ (.B1(net963),
    .Y(_04711_),
    .A1(net971),
    .A2(_04710_));
 sg13g2_nor3_1 _10706_ (.A(_00368_),
    .B(net1027),
    .C(net1013),
    .Y(_04712_));
 sg13g2_a21oi_1 _10707_ (.A1(net926),
    .A2(_04711_),
    .Y(_04713_),
    .B1(_04712_));
 sg13g2_mux4_1 _10708_ (.S0(net1132),
    .A0(_00372_),
    .A1(_00374_),
    .A2(_00373_),
    .A3(_00375_),
    .S1(net1208),
    .X(_04714_));
 sg13g2_mux4_1 _10709_ (.S0(net1132),
    .A0(_00380_),
    .A1(_00382_),
    .A2(_00381_),
    .A3(_00383_),
    .S1(net1208),
    .X(_04715_));
 sg13g2_and2_1 _10710_ (.A(net969),
    .B(_04715_),
    .X(_04716_));
 sg13g2_nand2_1 _10711_ (.Y(_04717_),
    .A(net1128),
    .B(_00379_));
 sg13g2_nand2b_1 _10712_ (.Y(_04718_),
    .B(_00377_),
    .A_N(net1128));
 sg13g2_a21oi_1 _10713_ (.A1(_04717_),
    .A2(_04718_),
    .Y(_04719_),
    .B1(_04045_));
 sg13g2_nand2_1 _10714_ (.Y(_04720_),
    .A(net1128),
    .B(_00378_));
 sg13g2_nand2b_1 _10715_ (.Y(_04721_),
    .B(_00376_),
    .A_N(net1132));
 sg13g2_a22oi_1 _10716_ (.Y(_04722_),
    .B1(net1002),
    .B2(net1001),
    .A2(_04721_),
    .A1(_04720_));
 sg13g2_or4_1 _10717_ (.A(net945),
    .B(_04716_),
    .C(_04719_),
    .D(_04722_),
    .X(_04723_));
 sg13g2_a221oi_1 _10718_ (.B2(net966),
    .C1(_04723_),
    .B1(_04714_),
    .A1(_04709_),
    .Y(_04724_),
    .A2(_04713_));
 sg13g2_a21oi_2 _10719_ (.B1(_04724_),
    .Y(_04725_),
    .A2(_04705_),
    .A1(_04696_));
 sg13g2_buf_2 fanout709 (.A(net711),
    .X(net709));
 sg13g2_a22oi_1 _10721_ (.Y(_04727_),
    .B1(net878),
    .B2(net899),
    .A2(_03177_),
    .A1(_03049_));
 sg13g2_nand3_1 _10722_ (.B(_03177_),
    .C(_04634_),
    .A(_03049_),
    .Y(_04728_));
 sg13g2_o21ai_1 _10723_ (.B1(_04104_),
    .Y(_04729_),
    .A1(net1101),
    .A2(net931));
 sg13g2_buf_2 fanout708 (.A(_08512_),
    .X(net708));
 sg13g2_nand2_1 _10725_ (.Y(_04731_),
    .A(net899),
    .B(_04729_));
 sg13g2_or2_1 _10726_ (.X(_04732_),
    .B(_04729_),
    .A(net904));
 sg13g2_mux2_1 _10727_ (.A0(_04731_),
    .A1(_04732_),
    .S(net872),
    .X(_04733_));
 sg13g2_nand3b_1 _10728_ (.B(_04728_),
    .C(_04733_),
    .Y(_04734_),
    .A_N(_04727_));
 sg13g2_buf_1 fanout707 (.A(net708),
    .X(net707));
 sg13g2_nand2_2 _10730_ (.Y(_04736_),
    .A(_04725_),
    .B(_04734_));
 sg13g2_buf_2 fanout706 (.A(net707),
    .X(net706));
 sg13g2_or2_1 _10732_ (.X(_04738_),
    .B(_04734_),
    .A(_04725_));
 sg13g2_buf_2 fanout705 (.A(net708),
    .X(net705));
 sg13g2_or2_1 _10734_ (.X(_04740_),
    .B(_00384_),
    .A(net1150));
 sg13g2_nor2b_1 _10735_ (.A(_00386_),
    .B_N(net1150),
    .Y(_04741_));
 sg13g2_o21ai_1 _10736_ (.B1(_04741_),
    .Y(_04742_),
    .A1(net1030),
    .A2(net1016));
 sg13g2_a21o_1 _10737_ (.A2(_04742_),
    .A1(_04740_),
    .B1(net1216),
    .X(_04743_));
 sg13g2_mux2_1 _10738_ (.A0(_00385_),
    .A1(_00387_),
    .S(net1152),
    .X(_04744_));
 sg13g2_o21ai_1 _10739_ (.B1(net964),
    .Y(_04745_),
    .A1(net974),
    .A2(_04744_));
 sg13g2_nor3_1 _10740_ (.A(_00384_),
    .B(net1030),
    .C(net1016),
    .Y(_04746_));
 sg13g2_a21oi_1 _10741_ (.A1(net932),
    .A2(_04745_),
    .Y(_04747_),
    .B1(_04746_));
 sg13g2_mux4_1 _10742_ (.S0(net1150),
    .A0(_00388_),
    .A1(_00390_),
    .A2(_00389_),
    .A3(_00391_),
    .S1(net1216),
    .X(_04748_));
 sg13g2_inv_1 _10743_ (.Y(_04749_),
    .A(_04748_));
 sg13g2_mux4_1 _10744_ (.S0(net1150),
    .A0(_00392_),
    .A1(_00394_),
    .A2(_00393_),
    .A3(_00395_),
    .S1(net1218),
    .X(_04750_));
 sg13g2_nand2_1 _10745_ (.Y(_04751_),
    .A(net991),
    .B(_04750_));
 sg13g2_o21ai_1 _10746_ (.B1(_04751_),
    .Y(_04752_),
    .A1(_04115_),
    .A2(_04749_));
 sg13g2_mux2_1 _10747_ (.A0(_00396_),
    .A1(_00398_),
    .S(net1152),
    .X(_04753_));
 sg13g2_nand3_1 _10748_ (.B(_03935_),
    .C(_04753_),
    .A(net1398),
    .Y(_04754_));
 sg13g2_mux2_1 _10749_ (.A0(_00397_),
    .A1(_00399_),
    .S(net1152),
    .X(_04755_));
 sg13g2_nand2b_1 _10750_ (.Y(_04756_),
    .B(_04755_),
    .A_N(_03711_));
 sg13g2_nand4_1 _10751_ (.B(_04009_),
    .C(_04754_),
    .A(net932),
    .Y(_04757_),
    .D(_04756_));
 sg13g2_a22oi_1 _10752_ (.Y(_04758_),
    .B1(_04752_),
    .B2(_04757_),
    .A2(_04747_),
    .A1(_04743_));
 sg13g2_buf_2 fanout704 (.A(net708),
    .X(net704));
 sg13g2_or2_1 _10754_ (.X(_04760_),
    .B(_00400_),
    .A(net1154));
 sg13g2_nor2b_1 _10755_ (.A(_00402_),
    .B_N(net1154),
    .Y(_04761_));
 sg13g2_o21ai_1 _10756_ (.B1(_04761_),
    .Y(_04762_),
    .A1(net1026),
    .A2(net1012));
 sg13g2_a21o_1 _10757_ (.A2(_04762_),
    .A1(_04760_),
    .B1(net1217),
    .X(_04763_));
 sg13g2_mux2_1 _10758_ (.A0(_00401_),
    .A1(_00403_),
    .S(net1154),
    .X(_04764_));
 sg13g2_o21ai_1 _10759_ (.B1(net964),
    .Y(_04765_),
    .A1(net974),
    .A2(_04764_));
 sg13g2_nor3_1 _10760_ (.A(_00400_),
    .B(net1031),
    .C(net1017),
    .Y(_04766_));
 sg13g2_a21oi_1 _10761_ (.A1(net932),
    .A2(_04765_),
    .Y(_04767_),
    .B1(_04766_));
 sg13g2_mux4_1 _10762_ (.S0(net1160),
    .A0(_00412_),
    .A1(_00414_),
    .A2(_00413_),
    .A3(_00415_),
    .S1(net1222),
    .X(_04768_));
 sg13g2_nand2_1 _10763_ (.Y(_04769_),
    .A(net1154),
    .B(_00407_));
 sg13g2_nand2b_1 _10764_ (.Y(_04770_),
    .B(_00405_),
    .A_N(net1154));
 sg13g2_a22oi_1 _10765_ (.Y(_04771_),
    .B1(net970),
    .B2(_03735_),
    .A2(_04770_),
    .A1(_04769_));
 sg13g2_nand2_1 _10766_ (.Y(_04772_),
    .A(net1134),
    .B(_00406_));
 sg13g2_nand2b_1 _10767_ (.Y(_04773_),
    .B(_00404_),
    .A_N(net1134));
 sg13g2_a22oi_1 _10768_ (.Y(_04774_),
    .B1(net1209),
    .B2(_03735_),
    .A2(_04773_),
    .A1(_04772_));
 sg13g2_mux4_1 _10769_ (.S0(net1153),
    .A0(_00408_),
    .A1(_00410_),
    .A2(_00409_),
    .A3(_00411_),
    .S1(net1217),
    .X(_04775_));
 sg13g2_and2_1 _10770_ (.A(net991),
    .B(_04775_),
    .X(_04776_));
 sg13g2_or4_1 _10771_ (.A(net946),
    .B(_04771_),
    .C(_04774_),
    .D(_04776_),
    .X(_04777_));
 sg13g2_a221oi_1 _10772_ (.B2(net969),
    .C1(_04777_),
    .B1(_04768_),
    .A1(_04763_),
    .Y(_04778_),
    .A2(_04767_));
 sg13g2_buf_2 fanout703 (.A(net708),
    .X(net703));
 sg13g2_nor2_1 _10774_ (.A(_04758_),
    .B(_04778_),
    .Y(_04780_));
 sg13g2_buf_2 fanout702 (.A(net703),
    .X(net702));
 sg13g2_nor2_1 _10776_ (.A(net949),
    .B(_03155_),
    .Y(_04782_));
 sg13g2_or3_1 _10777_ (.A(net949),
    .B(_03155_),
    .C(net899),
    .X(_04783_));
 sg13g2_a21oi_1 _10778_ (.A1(net899),
    .A2(_03895_),
    .Y(_04784_),
    .B1(net879));
 sg13g2_nor3_1 _10779_ (.A(net872),
    .B(net904),
    .C(_04052_),
    .Y(_04785_));
 sg13g2_a221oi_1 _10780_ (.B2(_04784_),
    .C1(_04785_),
    .B1(_04783_),
    .A1(_04634_),
    .Y(_04786_),
    .A2(_04782_));
 sg13g2_buf_1 fanout701 (.A(net702),
    .X(net701));
 sg13g2_xnor2_1 _10782_ (.Y(_04788_),
    .A(net620),
    .B(_04786_));
 sg13g2_nand3_1 _10783_ (.B(_04738_),
    .C(_04788_),
    .A(_04736_),
    .Y(_04789_));
 sg13g2_nor4_1 _10784_ (.A(_04600_),
    .B(_04642_),
    .C(_04690_),
    .D(_04789_),
    .Y(_04790_));
 sg13g2_nor2_2 _10785_ (.A(net1399),
    .B(net945),
    .Y(_04791_));
 sg13g2_nor2b_1 _10786_ (.A(net1167),
    .B_N(_00562_),
    .Y(_04792_));
 sg13g2_a22oi_1 _10787_ (.Y(_04793_),
    .B1(net1008),
    .B2(_04792_),
    .A2(_00564_),
    .A1(net1167));
 sg13g2_nor2b_1 _10788_ (.A(net1179),
    .B_N(_00563_),
    .Y(_04794_));
 sg13g2_a22oi_1 _10789_ (.Y(_04795_),
    .B1(_03683_),
    .B2(_04794_),
    .A2(_00565_),
    .A1(net1167));
 sg13g2_nor2b_1 _10790_ (.A(net1167),
    .B_N(_00558_),
    .Y(_04796_));
 sg13g2_a22oi_1 _10791_ (.Y(_04797_),
    .B1(net999),
    .B2(_04796_),
    .A2(_00560_),
    .A1(net1167));
 sg13g2_nor2b_1 _10792_ (.A(net1167),
    .B_N(_00559_),
    .Y(_04798_));
 sg13g2_a22oi_1 _10793_ (.Y(_04799_),
    .B1(net1005),
    .B2(_04798_),
    .A2(_00561_),
    .A1(net1167));
 sg13g2_nor4_1 _10794_ (.A(_04793_),
    .B(_04795_),
    .C(_04797_),
    .D(_04799_),
    .Y(_04800_));
 sg13g2_mux4_1 _10795_ (.S0(net1179),
    .A0(_00554_),
    .A1(_00556_),
    .A2(_00555_),
    .A3(_00557_),
    .S1(net1227),
    .X(_04801_));
 sg13g2_mux4_1 _10796_ (.S0(net1178),
    .A0(_00550_),
    .A1(_00552_),
    .A2(_00551_),
    .A3(_00553_),
    .S1(net1227),
    .X(_04802_));
 sg13g2_mux2_1 _10797_ (.A0(_04801_),
    .A1(_04802_),
    .S(net962),
    .X(_04803_));
 sg13g2_nor2_1 _10798_ (.A(net1394),
    .B(_03925_),
    .Y(_04804_));
 sg13g2_mux4_1 _10799_ (.S0(net1178),
    .A0(_00546_),
    .A1(_00548_),
    .A2(_00547_),
    .A3(_00549_),
    .S1(net1227),
    .X(_04805_));
 sg13g2_nand3_1 _10800_ (.B(net968),
    .C(_04805_),
    .A(net996),
    .Y(_04806_));
 sg13g2_nor3_1 _10801_ (.A(_00542_),
    .B(net1034),
    .C(net1020),
    .Y(_04807_));
 sg13g2_a21oi_1 _10802_ (.A1(net935),
    .A2(_04806_),
    .Y(_04808_),
    .B1(_04807_));
 sg13g2_a221oi_1 _10803_ (.B2(_04804_),
    .C1(_04808_),
    .B1(_04803_),
    .A1(_04791_),
    .Y(_04809_),
    .A2(_04800_));
 sg13g2_buf_2 fanout700 (.A(net702),
    .X(net700));
 sg13g2_mux4_1 _10805_ (.S0(net1179),
    .A0(_00567_),
    .A1(_00569_),
    .A2(_00571_),
    .A3(_00573_),
    .S1(net1114),
    .X(_04811_));
 sg13g2_inv_1 _10806_ (.Y(_04812_),
    .A(_04811_));
 sg13g2_nor2b_1 _10807_ (.A(net1179),
    .B_N(_00570_),
    .Y(_04813_));
 sg13g2_a22oi_1 _10808_ (.Y(_04814_),
    .B1(net1008),
    .B2(_04813_),
    .A2(_00572_),
    .A1(net1179));
 sg13g2_a22oi_1 _10809_ (.Y(_04815_),
    .B1(_04814_),
    .B2(net916),
    .A2(_04812_),
    .A1(net1227));
 sg13g2_or2_1 _10810_ (.X(_04816_),
    .B(_00566_),
    .A(net1168));
 sg13g2_nor2b_1 _10811_ (.A(_00568_),
    .B_N(net1168),
    .Y(_04817_));
 sg13g2_o21ai_1 _10812_ (.B1(_04817_),
    .Y(_04818_),
    .A1(net1034),
    .A2(net1020));
 sg13g2_a21o_1 _10813_ (.A2(_04818_),
    .A1(_04816_),
    .B1(net999),
    .X(_04819_));
 sg13g2_a21o_1 _10814_ (.A2(_00544_),
    .A1(net1178),
    .B1(net1227),
    .X(_04820_));
 sg13g2_o21ai_1 _10815_ (.B1(_04820_),
    .Y(_04821_),
    .A1(net1034),
    .A2(net1020));
 sg13g2_nand2_1 _10816_ (.Y(_04822_),
    .A(net959),
    .B(_00542_));
 sg13g2_nand2_2 _10817_ (.Y(_04823_),
    .A(net995),
    .B(net965));
 sg13g2_nor2b_1 _10818_ (.A(net1169),
    .B_N(_00543_),
    .Y(_04824_));
 sg13g2_a22oi_1 _10819_ (.Y(_04825_),
    .B1(_04824_),
    .B2(net976),
    .A2(_00545_),
    .A1(net1169));
 sg13g2_a22oi_1 _10820_ (.Y(_04826_),
    .B1(_04823_),
    .B2(_04825_),
    .A2(_04822_),
    .A1(_04821_));
 sg13g2_nand2_1 _10821_ (.Y(_04827_),
    .A(net939),
    .B(_03746_));
 sg13g2_buf_1 fanout699 (.A(_02111_),
    .X(net699));
 sg13g2_a22oi_1 _10823_ (.Y(_04829_),
    .B1(_04826_),
    .B2(net895),
    .A2(_04819_),
    .A1(_04815_));
 sg13g2_nand2_2 _10824_ (.Y(_04830_),
    .A(_04809_),
    .B(_04829_));
 sg13g2_buf_1 fanout698 (.A(net699),
    .X(net698));
 sg13g2_nand4_1 _10826_ (.B(_02955_),
    .C(_02964_),
    .A(_02951_),
    .Y(_04832_),
    .D(_02973_));
 sg13g2_buf_2 fanout697 (.A(net698),
    .X(net697));
 sg13g2_a21o_1 _10828_ (.A2(net896),
    .A1(net1235),
    .B1(net898),
    .X(_04834_));
 sg13g2_buf_2 fanout696 (.A(net699),
    .X(net696));
 sg13g2_mux2_1 _10830_ (.A0(_04832_),
    .A1(_04834_),
    .S(net901),
    .X(_04836_));
 sg13g2_xnor2_1 _10831_ (.Y(_04837_),
    .A(net876),
    .B(_04836_));
 sg13g2_xnor2_1 _10832_ (.Y(_04838_),
    .A(_04830_),
    .B(_04837_));
 sg13g2_a21oi_2 _10833_ (.B1(net897),
    .Y(_04839_),
    .A2(_04488_),
    .A1(net1238));
 sg13g2_mux2_1 _10834_ (.A0(_02946_),
    .A1(_04839_),
    .S(net901),
    .X(_04840_));
 sg13g2_xnor2_1 _10835_ (.Y(_04841_),
    .A(net876),
    .B(_04840_));
 sg13g2_nor2_1 _10836_ (.A(net1143),
    .B(_00598_),
    .Y(_04842_));
 sg13g2_nor3_1 _10837_ (.A(net958),
    .B(_00600_),
    .C(net920),
    .Y(_04843_));
 sg13g2_o21ai_1 _10838_ (.B1(net1040),
    .Y(_04844_),
    .A1(_04842_),
    .A2(_04843_));
 sg13g2_mux4_1 _10839_ (.S0(net1146),
    .A0(_00599_),
    .A1(_00601_),
    .A2(_00603_),
    .A3(_00605_),
    .S1(net1108),
    .X(_04845_));
 sg13g2_nor2_1 _10840_ (.A(net972),
    .B(_04845_),
    .Y(_04846_));
 sg13g2_nor2b_1 _10841_ (.A(net1146),
    .B_N(_00602_),
    .Y(_04847_));
 sg13g2_a22oi_1 _10842_ (.Y(_04848_),
    .B1(net1009),
    .B2(_04847_),
    .A2(_00604_),
    .A1(net1146));
 sg13g2_nor3_1 _10843_ (.A(net917),
    .B(_04846_),
    .C(_04848_),
    .Y(_04849_));
 sg13g2_nand2_1 _10844_ (.Y(_04850_),
    .A(net1143),
    .B(_00593_));
 sg13g2_nand2b_1 _10845_ (.Y(_04851_),
    .B(_00591_),
    .A_N(net1143));
 sg13g2_nand3_1 _10846_ (.B(_04850_),
    .C(_04851_),
    .A(net1213),
    .Y(_04852_));
 sg13g2_nor3_1 _10847_ (.A(net1213),
    .B(net1148),
    .C(_00590_),
    .Y(_04853_));
 sg13g2_nor2_1 _10848_ (.A(net997),
    .B(_04853_),
    .Y(_04854_));
 sg13g2_nor3_1 _10849_ (.A(net1108),
    .B(net1397),
    .C(_04238_),
    .Y(_04855_));
 sg13g2_nand3_1 _10850_ (.B(_04854_),
    .C(_04855_),
    .A(_04852_),
    .Y(_04856_));
 sg13g2_nand2_1 _10851_ (.Y(_04857_),
    .A(net1144),
    .B(_00585_));
 sg13g2_nand2b_1 _10852_ (.Y(_04858_),
    .B(_00583_),
    .A_N(net1142));
 sg13g2_nand3_1 _10853_ (.B(_04857_),
    .C(_04858_),
    .A(net1213),
    .Y(_04859_));
 sg13g2_inv_1 _10854_ (.Y(_04860_),
    .A(_00582_));
 sg13g2_a21oi_1 _10855_ (.A1(_04860_),
    .A2(_03743_),
    .Y(_04861_),
    .B1(net1392));
 sg13g2_nor3_1 _10856_ (.A(net1108),
    .B(net1003),
    .C(_04238_),
    .Y(_04862_));
 sg13g2_nand3_1 _10857_ (.B(_04861_),
    .C(_04862_),
    .A(_04859_),
    .Y(_04863_));
 sg13g2_nand2_1 _10858_ (.Y(_04864_),
    .A(net1144),
    .B(_00577_));
 sg13g2_nand2b_1 _10859_ (.Y(_04865_),
    .B(_00575_),
    .A_N(net1146));
 sg13g2_a21oi_1 _10860_ (.A1(_04864_),
    .A2(_04865_),
    .Y(_04866_),
    .B1(net973));
 sg13g2_and2_1 _10861_ (.A(_00576_),
    .B(_04238_),
    .X(_04867_));
 sg13g2_o21ai_1 _10862_ (.B1(net994),
    .Y(_04868_),
    .A1(_04866_),
    .A2(_04867_));
 sg13g2_nand4_1 _10863_ (.B(net992),
    .C(_04859_),
    .A(_00584_),
    .Y(_04869_),
    .D(_04861_));
 sg13g2_nand4_1 _10864_ (.B(_04863_),
    .C(_04868_),
    .A(_04856_),
    .Y(_04870_),
    .D(_04869_));
 sg13g2_nor2b_1 _10865_ (.A(_04853_),
    .B_N(_00592_),
    .Y(_04871_));
 sg13g2_nand4_1 _10866_ (.B(net915),
    .C(_04852_),
    .A(net929),
    .Y(_04872_),
    .D(_04871_));
 sg13g2_nor2_1 _10867_ (.A(net1391),
    .B(_04143_),
    .Y(_04873_));
 sg13g2_mux4_1 _10868_ (.S0(net1148),
    .A0(_00586_),
    .A1(_00588_),
    .A2(_00587_),
    .A3(_00589_),
    .S1(net1213),
    .X(_04874_));
 sg13g2_nand2_1 _10869_ (.Y(_04875_),
    .A(_00575_),
    .B(_00574_));
 sg13g2_a22oi_1 _10870_ (.Y(_04876_),
    .B1(_04410_),
    .B2(net989),
    .A2(_04875_),
    .A1(net1214));
 sg13g2_a22oi_1 _10871_ (.Y(_04877_),
    .B1(_04876_),
    .B2(net920),
    .A2(_04874_),
    .A1(_04873_));
 sg13g2_mux4_1 _10872_ (.S0(net1143),
    .A0(_00594_),
    .A1(_00596_),
    .A2(_00595_),
    .A3(_00597_),
    .S1(net1213),
    .X(_04878_));
 sg13g2_mux4_1 _10873_ (.S0(net1142),
    .A0(_00578_),
    .A1(_00580_),
    .A2(_00579_),
    .A3(_00581_),
    .S1(net1213),
    .X(_04879_));
 sg13g2_mux2_1 _10874_ (.A0(_04878_),
    .A1(_04879_),
    .S(net995),
    .X(_04880_));
 sg13g2_nand2b_1 _10875_ (.Y(_04881_),
    .B(_04880_),
    .A_N(_04115_));
 sg13g2_nand3_1 _10876_ (.B(_04877_),
    .C(_04881_),
    .A(_04872_),
    .Y(_04882_));
 sg13g2_a221oi_1 _10877_ (.B2(net929),
    .C1(_04882_),
    .B1(_04870_),
    .A1(_04844_),
    .Y(_04883_),
    .A2(_04849_));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_xnor2_1 _10879_ (.Y(_04885_),
    .A(_04841_),
    .B(net618));
 sg13g2_nor2_1 _10880_ (.A(_04305_),
    .B(_00632_),
    .Y(_04886_));
 sg13g2_nor2_1 _10881_ (.A(net1161),
    .B(_00630_),
    .Y(_04887_));
 sg13g2_a21oi_1 _10882_ (.A1(net929),
    .A2(_04886_),
    .Y(_04888_),
    .B1(_04887_));
 sg13g2_mux4_1 _10883_ (.S0(net1161),
    .A0(_00634_),
    .A1(_00636_),
    .A2(_00635_),
    .A3(_00637_),
    .S1(net1223),
    .X(_04889_));
 sg13g2_inv_1 _10884_ (.Y(_04890_),
    .A(_04889_));
 sg13g2_nor2b_1 _10885_ (.A(net1190),
    .B_N(_00631_),
    .Y(_04891_));
 sg13g2_a22oi_1 _10886_ (.Y(_04892_),
    .B1(net1005),
    .B2(_04891_),
    .A2(_00633_),
    .A1(net1190));
 sg13g2_a22oi_1 _10887_ (.Y(_04893_),
    .B1(_04892_),
    .B2(net917),
    .A2(_04890_),
    .A1(net1110));
 sg13g2_o21ai_1 _10888_ (.B1(_04893_),
    .Y(_04894_),
    .A1(net1000),
    .A2(_04888_));
 sg13g2_nor2_1 _10889_ (.A(net959),
    .B(_00616_),
    .Y(_04895_));
 sg13g2_nor2_1 _10890_ (.A(net1172),
    .B(_00614_),
    .Y(_04896_));
 sg13g2_a21oi_1 _10891_ (.A1(net936),
    .A2(_04895_),
    .Y(_04897_),
    .B1(_04896_));
 sg13g2_mux4_1 _10892_ (.S0(net1173),
    .A0(_00615_),
    .A1(_00617_),
    .A2(_00619_),
    .A3(_00621_),
    .S1(net1112),
    .X(_04898_));
 sg13g2_inv_1 _10893_ (.Y(_04899_),
    .A(_04898_));
 sg13g2_nor2b_1 _10894_ (.A(net1173),
    .B_N(_00618_),
    .Y(_04900_));
 sg13g2_a22oi_1 _10895_ (.Y(_04901_),
    .B1(net1009),
    .B2(_04900_),
    .A2(_00620_),
    .A1(net1173));
 sg13g2_a22oi_1 _10896_ (.Y(_04902_),
    .B1(_04901_),
    .B2(net948),
    .A2(_04899_),
    .A1(net1226));
 sg13g2_o21ai_1 _10897_ (.B1(_04902_),
    .Y(_04903_),
    .A1(_03725_),
    .A2(_04897_));
 sg13g2_or2_1 _10898_ (.X(_04904_),
    .B(_00606_),
    .A(net1188));
 sg13g2_nor2b_1 _10899_ (.A(_00608_),
    .B_N(net1190),
    .Y(_04905_));
 sg13g2_o21ai_1 _10900_ (.B1(_04905_),
    .Y(_04906_),
    .A1(net1036),
    .A2(net1022));
 sg13g2_a21o_1 _10901_ (.A2(_04906_),
    .A1(_04904_),
    .B1(net1235),
    .X(_04907_));
 sg13g2_mux2_1 _10902_ (.A0(_00607_),
    .A1(_00609_),
    .S(net1188),
    .X(_04908_));
 sg13g2_o21ai_1 _10903_ (.B1(net994),
    .Y(_04909_),
    .A1(net980),
    .A2(_04908_));
 sg13g2_nor3_1 _10904_ (.A(_00606_),
    .B(net1036),
    .C(net1022),
    .Y(_04910_));
 sg13g2_a21oi_1 _10905_ (.A1(net939),
    .A2(_04909_),
    .Y(_04911_),
    .B1(_04910_));
 sg13g2_or2_1 _10906_ (.X(_04912_),
    .B(net1188),
    .A(net1235));
 sg13g2_nor2b_1 _10907_ (.A(net1122),
    .B_N(_00622_),
    .Y(_04913_));
 sg13g2_a22oi_1 _10908_ (.Y(_04914_),
    .B1(_04912_),
    .B2(_04913_),
    .A2(_00626_),
    .A1(net1122));
 sg13g2_nor2b_1 _10909_ (.A(net1111),
    .B_N(_00624_),
    .Y(_04915_));
 sg13g2_a22oi_1 _10910_ (.Y(_04916_),
    .B1(_04477_),
    .B2(_04915_),
    .A2(_00628_),
    .A1(net1122));
 sg13g2_nor2b_1 _10911_ (.A(net1122),
    .B_N(_00623_),
    .Y(_04917_));
 sg13g2_a22oi_1 _10912_ (.Y(_04918_),
    .B1(net990),
    .B2(_04917_),
    .A2(_00627_),
    .A1(net1122));
 sg13g2_nor2b_1 _10913_ (.A(net1122),
    .B_N(_00625_),
    .Y(_04919_));
 sg13g2_a22oi_1 _10914_ (.Y(_04920_),
    .B1(net987),
    .B2(_04919_),
    .A2(_00629_),
    .A1(net1122));
 sg13g2_nor4_1 _10915_ (.A(_04914_),
    .B(_04916_),
    .C(_04918_),
    .D(_04920_),
    .Y(_04921_));
 sg13g2_mux2_1 _10916_ (.A0(_00611_),
    .A1(_00613_),
    .S(net1190),
    .X(_04922_));
 sg13g2_nand4_1 _10917_ (.B(net997),
    .C(net968),
    .A(net1235),
    .Y(_04923_),
    .D(_04922_));
 sg13g2_mux2_1 _10918_ (.A0(_00610_),
    .A1(_00612_),
    .S(net1188),
    .X(_04924_));
 sg13g2_nand3_1 _10919_ (.B(_04577_),
    .C(_04924_),
    .A(_03935_),
    .Y(_04925_));
 sg13g2_nand4_1 _10920_ (.B(_03746_),
    .C(_04923_),
    .A(net936),
    .Y(_04926_),
    .D(_04925_));
 sg13g2_a221oi_1 _10921_ (.B2(_04791_),
    .C1(_04926_),
    .B1(_04921_),
    .A1(_04907_),
    .Y(_04927_),
    .A2(_04911_));
 sg13g2_and3_2 _10922_ (.X(_04928_),
    .A(_04894_),
    .B(_04903_),
    .C(_04927_));
 sg13g2_buf_2 fanout694 (.A(net699),
    .X(net694));
 sg13g2_nor4_1 _10924_ (.A(_02882_),
    .B(_02888_),
    .C(_02897_),
    .D(net902),
    .Y(_04930_));
 sg13g2_a22oi_1 _10925_ (.Y(_04931_),
    .B1(net898),
    .B2(net911),
    .A2(net896),
    .A1(net1240));
 sg13g2_a21oi_1 _10926_ (.A1(_02916_),
    .A2(_04930_),
    .Y(_04932_),
    .B1(_04931_));
 sg13g2_xnor2_1 _10927_ (.Y(_04933_),
    .A(net882),
    .B(_04932_));
 sg13g2_xnor2_1 _10928_ (.Y(_04934_),
    .A(_04928_),
    .B(_04933_));
 sg13g2_buf_2 fanout693 (.A(net694),
    .X(net693));
 sg13g2_nor2b_1 _10930_ (.A(_00664_),
    .B_N(net1185),
    .Y(_04936_));
 sg13g2_o21ai_1 _10931_ (.B1(_04936_),
    .Y(_04937_),
    .A1(net1038),
    .A2(net1023));
 sg13g2_o21ai_1 _10932_ (.B1(_04937_),
    .Y(_04938_),
    .A1(net1185),
    .A2(_00662_));
 sg13g2_mux2_1 _10933_ (.A0(_00663_),
    .A1(_00665_),
    .S(net1187),
    .X(_04939_));
 sg13g2_mux4_1 _10934_ (.S0(net1186),
    .A0(_00666_),
    .A1(_00668_),
    .A2(_00667_),
    .A3(_00669_),
    .S1(net1229),
    .X(_04940_));
 sg13g2_nand2b_1 _10935_ (.Y(_04941_),
    .B(net1115),
    .A_N(_04940_));
 sg13g2_o21ai_1 _10936_ (.B1(_04941_),
    .Y(_04942_),
    .A1(net1005),
    .A2(_04939_));
 sg13g2_a22oi_1 _10937_ (.Y(_04943_),
    .B1(_04942_),
    .B2(net916),
    .A2(_04938_),
    .A1(net1041));
 sg13g2_mux4_1 _10938_ (.S0(net1187),
    .A0(_00654_),
    .A1(_00656_),
    .A2(_00655_),
    .A3(_00657_),
    .S1(net1229),
    .X(_04944_));
 sg13g2_nand3_1 _10939_ (.B(net914),
    .C(_04944_),
    .A(net937),
    .Y(_04945_));
 sg13g2_mux4_1 _10940_ (.S0(net1185),
    .A0(_00658_),
    .A1(_00660_),
    .A2(_00659_),
    .A3(_00661_),
    .S1(net1230),
    .X(_04946_));
 sg13g2_nand3_1 _10941_ (.B(net925),
    .C(_04946_),
    .A(net937),
    .Y(_04947_));
 sg13g2_nand2_1 _10942_ (.Y(_04948_),
    .A(net1194),
    .B(_00645_));
 sg13g2_nand2b_1 _10943_ (.Y(_04949_),
    .B(_00643_),
    .A_N(net1194));
 sg13g2_a22oi_1 _10944_ (.Y(_04950_),
    .B1(net1006),
    .B2(net988),
    .A2(_04949_),
    .A1(_04948_));
 sg13g2_nand2_1 _10945_ (.Y(_04951_),
    .A(net1185),
    .B(_00644_));
 sg13g2_nand2b_1 _10946_ (.Y(_04952_),
    .B(_00642_),
    .A_N(net1194));
 sg13g2_a22oi_1 _10947_ (.Y(_04953_),
    .B1(net1009),
    .B2(net988),
    .A2(_04952_),
    .A1(_04951_));
 sg13g2_nor2_1 _10948_ (.A(_04950_),
    .B(_04953_),
    .Y(_04954_));
 sg13g2_nand4_1 _10949_ (.B(_04945_),
    .C(_04947_),
    .A(net912),
    .Y(_04955_),
    .D(_04954_));
 sg13g2_nor2b_1 _10950_ (.A(_00648_),
    .B_N(net1191),
    .Y(_04956_));
 sg13g2_o21ai_1 _10951_ (.B1(_04956_),
    .Y(_04957_),
    .A1(net1038),
    .A2(net1020));
 sg13g2_o21ai_1 _10952_ (.B1(_04957_),
    .Y(_04958_),
    .A1(net1191),
    .A2(_00646_));
 sg13g2_mux4_1 _10953_ (.S0(net1191),
    .A0(_00647_),
    .A1(_00649_),
    .A2(_00651_),
    .A3(_00653_),
    .S1(net1117),
    .X(_04959_));
 sg13g2_nor2_1 _10954_ (.A(net978),
    .B(_04959_),
    .Y(_04960_));
 sg13g2_or2_1 _10955_ (.X(_04961_),
    .B(_04960_),
    .A(net948));
 sg13g2_nor2b_1 _10956_ (.A(net1192),
    .B_N(_00650_),
    .Y(_04962_));
 sg13g2_a22oi_1 _10957_ (.Y(_04963_),
    .B1(_04518_),
    .B2(_04962_),
    .A2(_00652_),
    .A1(net1192));
 sg13g2_a22oi_1 _10958_ (.Y(_04964_),
    .B1(_04961_),
    .B2(_04963_),
    .A2(_04958_),
    .A1(net1041));
 sg13g2_nor2b_1 _10959_ (.A(_00640_),
    .B_N(net1191),
    .Y(_04965_));
 sg13g2_o21ai_1 _10960_ (.B1(_04965_),
    .Y(_04966_),
    .A1(net1036),
    .A2(net1022));
 sg13g2_o21ai_1 _10961_ (.B1(_04966_),
    .Y(_04967_),
    .A1(net1191),
    .A2(_00638_));
 sg13g2_mux2_1 _10962_ (.A0(_00639_),
    .A1(_00641_),
    .S(net1191),
    .X(_04968_));
 sg13g2_o21ai_1 _10963_ (.B1(_03745_),
    .Y(_04969_),
    .A1(net980),
    .A2(_04968_));
 sg13g2_nor2_1 _10964_ (.A(_00638_),
    .B(net938),
    .Y(_04970_));
 sg13g2_a221oi_1 _10965_ (.B2(net938),
    .C1(_04970_),
    .B1(_04969_),
    .A1(net978),
    .Y(_04971_),
    .A2(_04967_));
 sg13g2_nor4_1 _10966_ (.A(_04943_),
    .B(_04955_),
    .C(_04964_),
    .D(_04971_),
    .Y(_04972_));
 sg13g2_buf_1 fanout692 (.A(net693),
    .X(net692));
 sg13g2_a22oi_1 _10968_ (.Y(_04974_),
    .B1(_02874_),
    .B2(net902),
    .A2(_02863_),
    .A1(_02855_));
 sg13g2_a22oi_1 _10969_ (.Y(_04975_),
    .B1(net898),
    .B2(net911),
    .A2(_04488_),
    .A1(net1242));
 sg13g2_a21oi_2 _10970_ (.B1(_04975_),
    .Y(_04976_),
    .A2(_04974_),
    .A1(_02848_));
 sg13g2_xnor2_1 _10971_ (.Y(_04977_),
    .A(net881),
    .B(_04976_));
 sg13g2_buf_2 fanout691 (.A(net693),
    .X(net691));
 sg13g2_xnor2_1 _10973_ (.Y(_04979_),
    .A(net615),
    .B(net403));
 sg13g2_and4_1 _10974_ (.A(_04838_),
    .B(_04885_),
    .C(_04934_),
    .D(_04979_),
    .X(_04980_));
 sg13g2_buf_2 fanout690 (.A(_02122_),
    .X(net690));
 sg13g2_nor2_2 _10976_ (.A(_04391_),
    .B(net919),
    .Y(_04982_));
 sg13g2_buf_2 fanout689 (.A(_02212_),
    .X(net689));
 sg13g2_mux2_1 _10978_ (.A0(_02781_),
    .A1(_04982_),
    .S(net901),
    .X(_04984_));
 sg13g2_xnor2_1 _10979_ (.Y(_04985_),
    .A(net876),
    .B(_04984_));
 sg13g2_inv_1 _10980_ (.Y(_04986_),
    .A(_04985_));
 sg13g2_nand2_1 _10981_ (.Y(_04987_),
    .A(net22),
    .B(net940));
 sg13g2_and2_1 _10982_ (.A(net901),
    .B(_04987_),
    .X(_04988_));
 sg13g2_a21oi_1 _10983_ (.A1(_02729_),
    .A2(net909),
    .Y(_04989_),
    .B1(_04988_));
 sg13g2_xnor2_1 _10984_ (.Y(_04990_),
    .A(net875),
    .B(_04989_));
 sg13g2_buf_2 fanout688 (.A(net689),
    .X(net688));
 sg13g2_mux4_1 _10986_ (.S0(net1188),
    .A0(_00791_),
    .A1(_00793_),
    .A2(_00795_),
    .A3(_00797_),
    .S1(net1122),
    .X(_04992_));
 sg13g2_nor2_1 _10987_ (.A(net980),
    .B(_04992_),
    .Y(_04993_));
 sg13g2_nor2b_1 _10988_ (.A(net1189),
    .B_N(_00794_),
    .Y(_04994_));
 sg13g2_a22oi_1 _10989_ (.Y(_04995_),
    .B1(net1009),
    .B2(_04994_),
    .A2(_00796_),
    .A1(net1189));
 sg13g2_inv_1 _10990_ (.Y(_04996_),
    .A(_00792_));
 sg13g2_o21ai_1 _10991_ (.B1(_04996_),
    .Y(_04997_),
    .A1(net1036),
    .A2(net1022));
 sg13g2_nor2b_1 _10992_ (.A(net1189),
    .B_N(_00790_),
    .Y(_04998_));
 sg13g2_a22oi_1 _10993_ (.Y(_04999_),
    .B1(_04998_),
    .B2(_03725_),
    .A2(_04997_),
    .A1(net1189));
 sg13g2_nor4_1 _10994_ (.A(net917),
    .B(_04993_),
    .C(_04995_),
    .D(_04999_),
    .Y(_05000_));
 sg13g2_nor3_1 _10995_ (.A(_00776_),
    .B(net921),
    .C(_03790_),
    .Y(_05001_));
 sg13g2_nor2b_1 _10996_ (.A(net1184),
    .B_N(_00778_),
    .Y(_05002_));
 sg13g2_a22oi_1 _10997_ (.Y(_05003_),
    .B1(_04518_),
    .B2(_05002_),
    .A2(_00780_),
    .A1(net1184));
 sg13g2_nor2_1 _10998_ (.A(_00774_),
    .B(_03781_),
    .Y(_05004_));
 sg13g2_nor2b_1 _10999_ (.A(net1112),
    .B_N(_00775_),
    .Y(_05005_));
 sg13g2_a22oi_1 _11000_ (.Y(_05006_),
    .B1(_03767_),
    .B2(_05005_),
    .A2(_00779_),
    .A1(net1112));
 sg13g2_nor2b_1 _11001_ (.A(net1112),
    .B_N(_00777_),
    .Y(_05007_));
 sg13g2_a22oi_1 _11002_ (.Y(_05008_),
    .B1(_03775_),
    .B2(_05007_),
    .A2(_00781_),
    .A1(net1113));
 sg13g2_or4_1 _11003_ (.A(net1003),
    .B(_05004_),
    .C(_05006_),
    .D(_05008_),
    .X(_05009_));
 sg13g2_nor4_2 _11004_ (.A(_03951_),
    .B(_05001_),
    .C(_05003_),
    .Y(_05010_),
    .D(_05009_));
 sg13g2_mux4_1 _11005_ (.S0(net1188),
    .A0(_00782_),
    .A1(_00784_),
    .A2(_00783_),
    .A3(_00785_),
    .S1(net1235),
    .X(_05011_));
 sg13g2_and3_1 _11006_ (.X(_05012_),
    .A(net939),
    .B(net914),
    .C(_05011_));
 sg13g2_mux4_1 _11007_ (.S0(net1188),
    .A0(_00786_),
    .A1(_00788_),
    .A2(_00787_),
    .A3(_00789_),
    .S1(net1235),
    .X(_05013_));
 sg13g2_and3_1 _11008_ (.X(_05014_),
    .A(net935),
    .B(net925),
    .C(_05013_));
 sg13g2_mux2_1 _11009_ (.A0(_00771_),
    .A1(_00773_),
    .S(net1188),
    .X(_05015_));
 sg13g2_nand4_1 _11010_ (.B(net997),
    .C(net968),
    .A(net1235),
    .Y(_05016_),
    .D(_05015_));
 sg13g2_mux2_1 _11011_ (.A0(_00770_),
    .A1(_00772_),
    .S(net1189),
    .X(_05017_));
 sg13g2_nand3_1 _11012_ (.B(_04577_),
    .C(_05017_),
    .A(_03935_),
    .Y(_05018_));
 sg13g2_nand4_1 _11013_ (.B(_03746_),
    .C(_05016_),
    .A(net939),
    .Y(_05019_),
    .D(_05018_));
 sg13g2_nor2_1 _11014_ (.A(_00768_),
    .B(_04477_),
    .Y(_05020_));
 sg13g2_nor2b_1 _11015_ (.A(net1176),
    .B_N(_00767_),
    .Y(_05021_));
 sg13g2_a22oi_1 _11016_ (.Y(_05022_),
    .B1(_05021_),
    .B2(net976),
    .A2(_00769_),
    .A1(net1176));
 sg13g2_o21ai_1 _11017_ (.B1(_03745_),
    .Y(_05023_),
    .A1(_00766_),
    .A2(_04912_));
 sg13g2_a22oi_1 _11018_ (.Y(_05024_),
    .B1(_05022_),
    .B2(_05023_),
    .A2(_05020_),
    .A1(net936));
 sg13g2_or4_1 _11019_ (.A(_05012_),
    .B(_05014_),
    .C(_05019_),
    .D(_05024_),
    .X(_05025_));
 sg13g2_or3_1 _11020_ (.A(_05000_),
    .B(_05010_),
    .C(_05025_),
    .X(_05026_));
 sg13g2_buf_1 fanout687 (.A(_02212_),
    .X(net687));
 sg13g2_nand2_2 _11022_ (.Y(_05028_),
    .A(net21),
    .B(net940));
 sg13g2_and2_1 _11023_ (.A(net901),
    .B(_05028_),
    .X(_05029_));
 sg13g2_a22oi_1 _11024_ (.Y(_05030_),
    .B1(_05029_),
    .B2(net875),
    .A2(net909),
    .A1(_02670_));
 sg13g2_buf_1 fanout686 (.A(net687),
    .X(net686));
 sg13g2_nand4_1 _11026_ (.B(_02634_),
    .C(_02658_),
    .A(_02603_),
    .Y(_05032_),
    .D(_02669_));
 sg13g2_nor2_1 _11027_ (.A(net909),
    .B(_05028_),
    .Y(_05033_));
 sg13g2_a22oi_1 _11028_ (.Y(_05034_),
    .B1(_05033_),
    .B2(net881),
    .A2(net909),
    .A1(_05032_));
 sg13g2_buf_2 fanout685 (.A(net687),
    .X(net685));
 sg13g2_nor3_2 _11030_ (.A(net613),
    .B(_05030_),
    .C(_05034_),
    .Y(_05036_));
 sg13g2_buf_2 fanout684 (.A(net687),
    .X(net684));
 sg13g2_nor2b_1 _11032_ (.A(net1184),
    .B_N(_00714_),
    .Y(_05038_));
 sg13g2_a22oi_1 _11033_ (.Y(_05039_),
    .B1(net1010),
    .B2(_05038_),
    .A2(_00716_),
    .A1(net1184));
 sg13g2_nor2_1 _11034_ (.A(net947),
    .B(_05039_),
    .Y(_05040_));
 sg13g2_nor3_1 _11035_ (.A(_00712_),
    .B(net924),
    .C(_03790_),
    .Y(_05041_));
 sg13g2_nor2b_1 _11036_ (.A(net1115),
    .B_N(_00713_),
    .Y(_05042_));
 sg13g2_a22oi_1 _11037_ (.Y(_05043_),
    .B1(net987),
    .B2(_05042_),
    .A2(_00717_),
    .A1(net1115));
 sg13g2_nor2b_1 _11038_ (.A(net1115),
    .B_N(_00711_),
    .Y(_05044_));
 sg13g2_a22oi_1 _11039_ (.Y(_05045_),
    .B1(net990),
    .B2(_05044_),
    .A2(_00715_),
    .A1(net1115));
 sg13g2_nor3_1 _11040_ (.A(net1229),
    .B(_00710_),
    .C(_04410_),
    .Y(_05046_));
 sg13g2_nor4_1 _11041_ (.A(_05041_),
    .B(_05043_),
    .C(_05045_),
    .D(_05046_),
    .Y(_05047_));
 sg13g2_nor2b_1 _11042_ (.A(net1184),
    .B_N(_00703_),
    .Y(_05048_));
 sg13g2_a22oi_1 _11043_ (.Y(_05049_),
    .B1(net1005),
    .B2(_05048_),
    .A2(_00705_),
    .A1(net1184));
 sg13g2_nor2b_1 _11044_ (.A(net1185),
    .B_N(_00707_),
    .Y(_05050_));
 sg13g2_a22oi_1 _11045_ (.Y(_05051_),
    .B1(net1006),
    .B2(_05050_),
    .A2(_00709_),
    .A1(net1185));
 sg13g2_nor2b_1 _11046_ (.A(net1185),
    .B_N(_00706_),
    .Y(_05052_));
 sg13g2_a22oi_1 _11047_ (.Y(_05053_),
    .B1(net1008),
    .B2(_05052_),
    .A2(_00708_),
    .A1(net1185));
 sg13g2_or4_1 _11048_ (.A(net989),
    .B(_05049_),
    .C(_05051_),
    .D(_05053_),
    .X(_05054_));
 sg13g2_nor2b_1 _11049_ (.A(_00702_),
    .B_N(_03783_),
    .Y(_05055_));
 sg13g2_nor3_1 _11050_ (.A(_00704_),
    .B(net921),
    .C(_03790_),
    .Y(_05056_));
 sg13g2_a22oi_1 _11051_ (.Y(_05057_),
    .B1(_05055_),
    .B2(_05056_),
    .A2(_05054_),
    .A1(net938));
 sg13g2_a21oi_2 _11052_ (.B1(_05057_),
    .Y(_05058_),
    .A2(_05047_),
    .A1(_05040_));
 sg13g2_mux4_1 _11053_ (.S0(net1194),
    .A0(_00722_),
    .A1(_00724_),
    .A2(_00723_),
    .A3(_00725_),
    .S1(net1234),
    .X(_05059_));
 sg13g2_nand2_1 _11054_ (.Y(_05060_),
    .A(net925),
    .B(_05059_));
 sg13g2_nor2b_2 _11055_ (.A(net1196),
    .B_N(net1119),
    .Y(_05061_));
 sg13g2_buf_1 fanout683 (.A(_02212_),
    .X(net683));
 sg13g2_nand3_1 _11057_ (.B(net993),
    .C(_05061_),
    .A(_00730_),
    .Y(_05063_));
 sg13g2_nand3_1 _11058_ (.B(net1401),
    .C(net1394),
    .A(net1120),
    .Y(_05064_));
 sg13g2_buf_1 fanout682 (.A(net683),
    .X(net682));
 sg13g2_a21oi_1 _11060_ (.A1(net1194),
    .A2(_00732_),
    .Y(_05066_),
    .B1(net1234));
 sg13g2_or2_1 _11061_ (.X(_05067_),
    .B(_05066_),
    .A(_05064_));
 sg13g2_nor2b_1 _11062_ (.A(net1194),
    .B_N(_00731_),
    .Y(_05068_));
 sg13g2_a22oi_1 _11063_ (.Y(_05069_),
    .B1(_05068_),
    .B2(net978),
    .A2(_00733_),
    .A1(net1195));
 sg13g2_a21o_1 _11064_ (.A2(_05067_),
    .A1(_05063_),
    .B1(_05069_),
    .X(_05070_));
 sg13g2_mux4_1 _11065_ (.S0(net1186),
    .A0(_00718_),
    .A1(_00720_),
    .A2(_00719_),
    .A3(_00721_),
    .S1(net1230),
    .X(_05071_));
 sg13g2_nand2_1 _11066_ (.Y(_05072_),
    .A(net914),
    .B(_05071_));
 sg13g2_nor2_1 _11067_ (.A(net1196),
    .B(net1119),
    .Y(_05073_));
 sg13g2_nand3_1 _11068_ (.B(net993),
    .C(_05073_),
    .A(_00726_),
    .Y(_05074_));
 sg13g2_nand3b_1 _11069_ (.B(net1401),
    .C(net1394),
    .Y(_05075_),
    .A_N(net1120));
 sg13g2_buf_2 fanout681 (.A(net683),
    .X(net681));
 sg13g2_a21oi_1 _11071_ (.A1(net1195),
    .A2(_00728_),
    .Y(_05077_),
    .B1(net1234));
 sg13g2_or2_1 _11072_ (.X(_05078_),
    .B(_05077_),
    .A(_05075_));
 sg13g2_nor2b_1 _11073_ (.A(net1195),
    .B_N(_00727_),
    .Y(_05079_));
 sg13g2_a22oi_1 _11074_ (.Y(_05080_),
    .B1(_05079_),
    .B2(net978),
    .A2(_00729_),
    .A1(net1195));
 sg13g2_a21o_1 _11075_ (.A2(_05078_),
    .A1(_05074_),
    .B1(_05080_),
    .X(_05081_));
 sg13g2_nand4_1 _11076_ (.B(_05070_),
    .C(_05072_),
    .A(_05060_),
    .Y(_05082_),
    .D(_05081_));
 sg13g2_nand2_1 _11077_ (.Y(_05083_),
    .A(net941),
    .B(_05082_));
 sg13g2_and3_1 _11078_ (.X(_05084_),
    .A(_03747_),
    .B(_05058_),
    .C(_05083_));
 sg13g2_buf_2 fanout680 (.A(net683),
    .X(net680));
 sg13g2_nor3_1 _11080_ (.A(_04990_),
    .B(_05036_),
    .C(_05084_),
    .Y(_05086_));
 sg13g2_o21ai_1 _11081_ (.B1(net402),
    .Y(_05087_),
    .A1(_04990_),
    .A2(_05036_));
 sg13g2_o21ai_1 _11082_ (.B1(_05087_),
    .Y(_05088_),
    .A1(_04986_),
    .A2(_05086_));
 sg13g2_nand2_1 _11083_ (.Y(_05089_),
    .A(net402),
    .B(_04985_));
 sg13g2_mux4_1 _11084_ (.S0(net1169),
    .A0(_00762_),
    .A1(_00764_),
    .A2(_00763_),
    .A3(_00765_),
    .S1(net1226),
    .X(_05090_));
 sg13g2_mux4_1 _11085_ (.S0(net1164),
    .A0(_00754_),
    .A1(_00756_),
    .A2(_00755_),
    .A3(_00757_),
    .S1(net1225),
    .X(_05091_));
 sg13g2_mux4_1 _11086_ (.S0(net1164),
    .A0(_00758_),
    .A1(_00760_),
    .A2(_00759_),
    .A3(_00761_),
    .S1(net1225),
    .X(_05092_));
 sg13g2_mux4_1 _11087_ (.S0(net1168),
    .A0(_00750_),
    .A1(_00752_),
    .A2(_00751_),
    .A3(_00753_),
    .S1(net1226),
    .X(_05093_));
 sg13g2_mux4_1 _11088_ (.S0(net1003),
    .A0(_05090_),
    .A1(_05091_),
    .A2(_05092_),
    .A3(_05093_),
    .S1(net962),
    .X(_05094_));
 sg13g2_nand2b_1 _11089_ (.Y(_05095_),
    .B(_05094_),
    .A_N(net946));
 sg13g2_nor3_1 _11090_ (.A(net959),
    .B(_00744_),
    .C(net998),
    .Y(_05096_));
 sg13g2_nor3_1 _11091_ (.A(net1177),
    .B(_00742_),
    .C(net998),
    .Y(_05097_));
 sg13g2_a21oi_1 _11092_ (.A1(net935),
    .A2(_05096_),
    .Y(_05098_),
    .B1(_05097_));
 sg13g2_nor2b_1 _11093_ (.A(net1165),
    .B_N(_00746_),
    .Y(_05099_));
 sg13g2_a22oi_1 _11094_ (.Y(_05100_),
    .B1(net1007),
    .B2(_05099_),
    .A2(_00748_),
    .A1(net1166));
 sg13g2_mux4_1 _11095_ (.S0(net1166),
    .A0(_00743_),
    .A1(_00745_),
    .A2(_00747_),
    .A3(_00749_),
    .S1(net1113),
    .X(_05101_));
 sg13g2_nor2_1 _11096_ (.A(net976),
    .B(_05101_),
    .Y(_05102_));
 sg13g2_a22oi_1 _11097_ (.Y(_05103_),
    .B1(_05102_),
    .B2(net947),
    .A2(_05100_),
    .A1(net935));
 sg13g2_nand2_1 _11098_ (.Y(_05104_),
    .A(_05098_),
    .B(_05103_));
 sg13g2_or2_1 _11099_ (.X(_05105_),
    .B(_04240_),
    .A(_00740_));
 sg13g2_inv_1 _11100_ (.Y(_05106_),
    .A(_00738_));
 sg13g2_nand2_1 _11101_ (.Y(_05107_),
    .A(net996),
    .B(net968));
 sg13g2_nor2b_1 _11102_ (.A(net1175),
    .B_N(_00739_),
    .Y(_05108_));
 sg13g2_a22oi_1 _11103_ (.Y(_05109_),
    .B1(_05108_),
    .B2(net977),
    .A2(_00741_),
    .A1(net1175));
 sg13g2_a22oi_1 _11104_ (.Y(_05110_),
    .B1(_05107_),
    .B2(_05109_),
    .A2(_03743_),
    .A1(_05106_));
 sg13g2_inv_1 _11105_ (.Y(_05111_),
    .A(_00737_));
 sg13g2_buf_2 fanout679 (.A(net680),
    .X(net679));
 sg13g2_o21ai_1 _11107_ (.B1(net959),
    .Y(_05113_),
    .A1(net976),
    .A2(_00735_));
 sg13g2_o21ai_1 _11108_ (.B1(_05113_),
    .Y(_05114_),
    .A1(_05111_),
    .A2(net987));
 sg13g2_mux2_1 _11109_ (.A0(_00734_),
    .A1(_00736_),
    .S(net1175),
    .X(_05115_));
 sg13g2_nand3_1 _11110_ (.B(_04577_),
    .C(_05115_),
    .A(net1041),
    .Y(_05116_));
 sg13g2_nand2_1 _11111_ (.Y(_05117_),
    .A(net936),
    .B(_05116_));
 sg13g2_a221oi_1 _11112_ (.B2(net994),
    .C1(_05117_),
    .B1(_05114_),
    .A1(_05105_),
    .Y(_05118_),
    .A2(_05110_));
 sg13g2_buf_1 fanout678 (.A(_02250_),
    .X(net678));
 sg13g2_and3_2 _11114_ (.X(_05120_),
    .A(_05095_),
    .B(_05104_),
    .C(_05118_));
 sg13g2_buf_2 fanout677 (.A(net678),
    .X(net677));
 sg13g2_a21oi_1 _11116_ (.A1(_04990_),
    .A2(_05036_),
    .Y(_05122_),
    .B1(_05120_));
 sg13g2_nor2_1 _11117_ (.A(net921),
    .B(_05107_),
    .Y(_05123_));
 sg13g2_inv_1 _11118_ (.Y(_05124_),
    .A(_00676_));
 sg13g2_o21ai_1 _11119_ (.B1(_05124_),
    .Y(_05125_),
    .A1(net1037),
    .A2(net1022));
 sg13g2_mux4_1 _11120_ (.S0(net979),
    .A0(_00675_),
    .A1(_00674_),
    .A2(_00677_),
    .A3(_05125_),
    .S1(net1201),
    .X(_05126_));
 sg13g2_mux4_1 _11121_ (.S0(net1200),
    .A0(_00686_),
    .A1(_00688_),
    .A2(_00687_),
    .A3(_00689_),
    .S1(net1232),
    .X(_05127_));
 sg13g2_a221oi_1 _11122_ (.B2(net915),
    .C1(net895),
    .B1(_05127_),
    .A1(_05123_),
    .Y(_05128_),
    .A2(_05126_));
 sg13g2_buf_2 fanout676 (.A(_02250_),
    .X(net676));
 sg13g2_nor3_1 _11124_ (.A(net960),
    .B(_00680_),
    .C(net1000),
    .Y(_05130_));
 sg13g2_mux4_1 _11125_ (.S0(net1193),
    .A0(_00679_),
    .A1(_00681_),
    .A2(_00683_),
    .A3(_00685_),
    .S1(net1117),
    .X(_05131_));
 sg13g2_nor2_1 _11126_ (.A(net978),
    .B(_05131_),
    .Y(_05132_));
 sg13g2_nor3_1 _11127_ (.A(net1193),
    .B(_00678_),
    .C(net1000),
    .Y(_05133_));
 sg13g2_a22oi_1 _11128_ (.Y(_05134_),
    .B1(_05132_),
    .B2(_05133_),
    .A2(_05130_),
    .A1(net942));
 sg13g2_nand2b_1 _11129_ (.Y(_05135_),
    .B(net1201),
    .A_N(_00684_));
 sg13g2_o21ai_1 _11130_ (.B1(_05135_),
    .Y(_05136_),
    .A1(net1201),
    .A2(_00682_));
 sg13g2_nand2_1 _11131_ (.Y(_05137_),
    .A(net1401),
    .B(net997));
 sg13g2_a22oi_1 _11132_ (.Y(_05138_),
    .B1(net922),
    .B2(_05137_),
    .A2(_05136_),
    .A1(_03935_));
 sg13g2_and2_1 _11133_ (.A(_05134_),
    .B(_05138_),
    .X(_05139_));
 sg13g2_nor2b_1 _11134_ (.A(_00696_),
    .B_N(net1199),
    .Y(_05140_));
 sg13g2_o21ai_1 _11135_ (.B1(_05140_),
    .Y(_05141_),
    .A1(net1037),
    .A2(net1022));
 sg13g2_o21ai_1 _11136_ (.B1(_05141_),
    .Y(_05142_),
    .A1(net1198),
    .A2(_00694_));
 sg13g2_mux2_1 _11137_ (.A0(_00698_),
    .A1(_00700_),
    .S(net1196),
    .X(_05143_));
 sg13g2_mux4_1 _11138_ (.S0(net1196),
    .A0(_00695_),
    .A1(_00697_),
    .A2(_00699_),
    .A3(_00701_),
    .S1(net1120),
    .X(_05144_));
 sg13g2_nand2b_1 _11139_ (.Y(_05145_),
    .B(net1232),
    .A_N(_05144_));
 sg13g2_o21ai_1 _11140_ (.B1(_05145_),
    .Y(_05146_),
    .A1(net1009),
    .A2(_05143_));
 sg13g2_a22oi_1 _11141_ (.Y(_05147_),
    .B1(_05146_),
    .B2(net917),
    .A2(_05142_),
    .A1(net1041));
 sg13g2_mux2_1 _11142_ (.A0(_00671_),
    .A1(_00673_),
    .S(net1193),
    .X(_05148_));
 sg13g2_o21ai_1 _11143_ (.B1(net994),
    .Y(_05149_),
    .A1(net980),
    .A2(_05148_));
 sg13g2_nor2b_1 _11144_ (.A(_00672_),
    .B_N(net1193),
    .Y(_05150_));
 sg13g2_o21ai_1 _11145_ (.B1(_05150_),
    .Y(_05151_),
    .A1(net1037),
    .A2(net1023));
 sg13g2_o21ai_1 _11146_ (.B1(_05151_),
    .Y(_05152_),
    .A1(net1189),
    .A2(_00670_));
 sg13g2_nor2_1 _11147_ (.A(_00670_),
    .B(net939),
    .Y(_05153_));
 sg13g2_a221oi_1 _11148_ (.B2(net980),
    .C1(_05153_),
    .B1(_05152_),
    .A1(net939),
    .Y(_05154_),
    .A2(_05149_));
 sg13g2_nor2b_1 _11149_ (.A(_00692_),
    .B_N(net1200),
    .Y(_05155_));
 sg13g2_o21ai_1 _11150_ (.B1(_05155_),
    .Y(_05156_),
    .A1(net1036),
    .A2(net1022));
 sg13g2_o21ai_1 _11151_ (.B1(_05156_),
    .Y(_05157_),
    .A1(net1200),
    .A2(_00690_));
 sg13g2_nor2b_1 _11152_ (.A(net1200),
    .B_N(_00691_),
    .Y(_05158_));
 sg13g2_a22oi_1 _11153_ (.Y(_05159_),
    .B1(_05158_),
    .B2(net978),
    .A2(_00693_),
    .A1(net1200));
 sg13g2_nand2_1 _11154_ (.Y(_05160_),
    .A(net943),
    .B(_03737_));
 sg13g2_a22oi_1 _11155_ (.Y(_05161_),
    .B1(_05159_),
    .B2(_05160_),
    .A2(_05157_),
    .A1(net979));
 sg13g2_nor4_2 _11156_ (.A(_05139_),
    .B(_05147_),
    .C(_05154_),
    .Y(_05162_),
    .D(_05161_));
 sg13g2_and2_1 _11157_ (.A(_05128_),
    .B(_05162_),
    .X(_05163_));
 sg13g2_buf_2 fanout675 (.A(net676),
    .X(net675));
 sg13g2_nand3_1 _11159_ (.B(net1251),
    .C(net1254),
    .A(net1375),
    .Y(_05165_));
 sg13g2_nand2_1 _11160_ (.Y(_05166_),
    .A(net30),
    .B(_02570_));
 sg13g2_a22oi_1 _11161_ (.Y(_05167_),
    .B1(_03812_),
    .B2(_03814_),
    .A2(_05166_),
    .A1(_05165_));
 sg13g2_nor2_2 _11162_ (.A(_04104_),
    .B(_03837_),
    .Y(_05168_));
 sg13g2_nor3_1 _11163_ (.A(net908),
    .B(_05167_),
    .C(_05168_),
    .Y(_05169_));
 sg13g2_a21oi_1 _11164_ (.A1(_02820_),
    .A2(net908),
    .Y(_05170_),
    .B1(_05169_));
 sg13g2_xnor2_1 _11165_ (.Y(_05171_),
    .A(net875),
    .B(_05170_));
 sg13g2_nor2_1 _11166_ (.A(net401),
    .B(_05171_),
    .Y(_05172_));
 sg13g2_a21oi_1 _11167_ (.A1(_05089_),
    .A2(_05122_),
    .Y(_05173_),
    .B1(_05172_));
 sg13g2_and2_1 _11168_ (.A(net401),
    .B(_05171_),
    .X(_05174_));
 sg13g2_a21o_1 _11169_ (.A2(_05173_),
    .A1(_05088_),
    .B1(_05174_),
    .X(_05175_));
 sg13g2_buf_2 fanout674 (.A(_02250_),
    .X(net674));
 sg13g2_and2_2 _11171_ (.A(_04809_),
    .B(_04829_),
    .X(_05177_));
 sg13g2_buf_2 fanout673 (.A(net674),
    .X(net673));
 sg13g2_nand2_1 _11173_ (.Y(_05179_),
    .A(_05177_),
    .B(_04837_));
 sg13g2_inv_1 _11174_ (.Y(_05180_),
    .A(_04841_));
 sg13g2_buf_2 fanout672 (.A(net674),
    .X(net672));
 sg13g2_nor2_1 _11176_ (.A(_05180_),
    .B(net619),
    .Y(_05182_));
 sg13g2_and2_1 _11177_ (.A(net876),
    .B(_04976_),
    .X(_05183_));
 sg13g2_or2_1 _11178_ (.X(_05184_),
    .B(_04932_),
    .A(_04928_));
 sg13g2_nand3_1 _11179_ (.B(_04903_),
    .C(_04927_),
    .A(_04894_),
    .Y(_05185_));
 sg13g2_buf_1 fanout671 (.A(net672),
    .X(net671));
 sg13g2_a22oi_1 _11181_ (.Y(_05187_),
    .B1(_04976_),
    .B2(net876),
    .A2(_04932_),
    .A1(_05185_));
 sg13g2_a21o_1 _11182_ (.A2(_05184_),
    .A1(_05183_),
    .B1(_05187_),
    .X(_05188_));
 sg13g2_xnor2_1 _11183_ (.Y(_05189_),
    .A(net882),
    .B(_04836_));
 sg13g2_o21ai_1 _11184_ (.B1(_04841_),
    .Y(_05190_),
    .A1(_04830_),
    .A2(_05189_));
 sg13g2_a21o_1 _11185_ (.A2(_04837_),
    .A1(_05177_),
    .B1(net619),
    .X(_05191_));
 sg13g2_nor2_1 _11186_ (.A(_05185_),
    .B(_04933_),
    .Y(_05192_));
 sg13g2_a221oi_1 _11187_ (.B2(_05191_),
    .C1(_05192_),
    .B1(_05190_),
    .A1(net616),
    .Y(_05193_),
    .A2(_05188_));
 sg13g2_nand2_1 _11188_ (.Y(_05194_),
    .A(_04830_),
    .B(_05189_));
 sg13g2_inv_1 _11189_ (.Y(_05195_),
    .A(_05194_));
 sg13g2_a22oi_1 _11190_ (.Y(_05196_),
    .B1(_05193_),
    .B2(_05195_),
    .A2(_05182_),
    .A1(_05179_));
 sg13g2_a21o_1 _11191_ (.A2(_05175_),
    .A1(_04980_),
    .B1(_05196_),
    .X(_05197_));
 sg13g2_a21oi_2 _11192_ (.B1(_04426_),
    .Y(_05198_),
    .A2(_04414_),
    .A1(_04405_));
 sg13g2_buf_2 fanout670 (.A(net671),
    .X(net670));
 sg13g2_nand2_2 _11194_ (.Y(_05200_),
    .A(_05198_),
    .B(_04442_));
 sg13g2_nor2_2 _11195_ (.A(_05198_),
    .B(_04442_),
    .Y(_05201_));
 sg13g2_a22oi_1 _11196_ (.Y(_05202_),
    .B1(_05201_),
    .B2(_04497_),
    .A2(_05200_),
    .A1(_04552_));
 sg13g2_nor3_1 _11197_ (.A(_04563_),
    .B(_04582_),
    .C(_04591_),
    .Y(_05203_));
 sg13g2_buf_2 fanout669 (.A(_02290_),
    .X(net669));
 sg13g2_and2_1 _11199_ (.A(_05203_),
    .B(_04597_),
    .X(_05205_));
 sg13g2_nand3_1 _11200_ (.B(_04500_),
    .C(_04501_),
    .A(_04502_),
    .Y(_05206_));
 sg13g2_buf_2 fanout668 (.A(net669),
    .X(net668));
 sg13g2_o21ai_1 _11202_ (.B1(_05206_),
    .Y(_05208_),
    .A1(_04503_),
    .A2(_05205_));
 sg13g2_inv_1 _11203_ (.Y(_05209_),
    .A(_04597_));
 sg13g2_o21ai_1 _11204_ (.B1(_05209_),
    .Y(_05210_),
    .A1(_04497_),
    .A2(net623));
 sg13g2_nand3b_1 _11205_ (.B(_05208_),
    .C(_05210_),
    .Y(_05211_),
    .A_N(_05202_));
 sg13g2_inv_1 _11206_ (.Y(_05212_),
    .A(_04786_));
 sg13g2_o21ai_1 _11207_ (.B1(_04738_),
    .Y(_05213_),
    .A1(_04780_),
    .A2(_05212_));
 sg13g2_a21oi_1 _11208_ (.A1(_05206_),
    .A2(_05209_),
    .Y(_05214_),
    .B1(net623));
 sg13g2_a21oi_2 _11209_ (.B1(_04684_),
    .Y(_05215_),
    .A2(_04662_),
    .A1(_04651_));
 sg13g2_buf_2 fanout667 (.A(_02294_),
    .X(net667));
 sg13g2_buf_1 fanout666 (.A(net667),
    .X(net666));
 sg13g2_nand3_1 _11212_ (.B(_04640_),
    .C(_04689_),
    .A(net621),
    .Y(_05218_));
 sg13g2_a21oi_1 _11213_ (.A1(net622),
    .A2(_04640_),
    .Y(_05219_),
    .B1(_04689_));
 sg13g2_a21oi_1 _11214_ (.A1(_05215_),
    .A2(_05218_),
    .Y(_05220_),
    .B1(_05219_));
 sg13g2_a22oi_1 _11215_ (.Y(_05221_),
    .B1(_05214_),
    .B2(_05220_),
    .A2(_05213_),
    .A1(_04736_));
 sg13g2_nor2_1 _11216_ (.A(_04642_),
    .B(_04690_),
    .Y(_05222_));
 sg13g2_a21o_2 _11217_ (.A2(_04705_),
    .A1(_04696_),
    .B1(_04724_),
    .X(_05223_));
 sg13g2_buf_2 fanout665 (.A(net666),
    .X(net665));
 sg13g2_or2_1 _11219_ (.X(_05225_),
    .B(_04778_),
    .A(_04758_));
 sg13g2_buf_2 fanout664 (.A(net667),
    .X(net664));
 sg13g2_nor3_1 _11221_ (.A(_05223_),
    .B(_05225_),
    .C(_04786_),
    .Y(_05227_));
 sg13g2_o21ai_1 _11222_ (.B1(_05223_),
    .Y(_05228_),
    .A1(_05225_),
    .A2(_04786_));
 sg13g2_o21ai_1 _11223_ (.B1(_05228_),
    .Y(_05229_),
    .A1(_04734_),
    .A2(_05227_));
 sg13g2_a21oi_1 _11224_ (.A1(_05222_),
    .A2(_05229_),
    .Y(_05230_),
    .B1(_05220_));
 sg13g2_a21oi_1 _11225_ (.A1(_05211_),
    .A2(_05221_),
    .Y(_05231_),
    .B1(_05230_));
 sg13g2_a21oi_1 _11226_ (.A1(_04790_),
    .A2(_05197_),
    .Y(_05232_),
    .B1(_05231_));
 sg13g2_xnor2_1 _11227_ (.Y(_05233_),
    .A(net402),
    .B(_04985_));
 sg13g2_xnor2_1 _11228_ (.Y(_05234_),
    .A(net401),
    .B(_05171_));
 sg13g2_buf_2 fanout663 (.A(net667),
    .X(net663));
 sg13g2_xnor2_1 _11230_ (.Y(_05236_),
    .A(_04990_),
    .B(_05120_));
 sg13g2_nor3_2 _11231_ (.A(_05000_),
    .B(_05010_),
    .C(_05025_),
    .Y(_05237_));
 sg13g2_buf_2 fanout662 (.A(net667),
    .X(net662));
 sg13g2_nor2_2 _11233_ (.A(_05030_),
    .B(_05034_),
    .Y(_05239_));
 sg13g2_buf_1 fanout661 (.A(net662),
    .X(net661));
 sg13g2_xnor2_1 _11235_ (.Y(_05241_),
    .A(_05237_),
    .B(_05239_));
 sg13g2_nor4_2 _11236_ (.A(_05233_),
    .B(_05234_),
    .C(_05236_),
    .Y(_05242_),
    .D(_05241_));
 sg13g2_and2_1 _11237_ (.A(_04980_),
    .B(_05242_),
    .X(_05243_));
 sg13g2_nor2_1 _11238_ (.A(net958),
    .B(_00920_),
    .Y(_05244_));
 sg13g2_nor2_1 _11239_ (.A(net1146),
    .B(_00918_),
    .Y(_05245_));
 sg13g2_a21oi_1 _11240_ (.A1(net929),
    .A2(_05244_),
    .Y(_05246_),
    .B1(_05245_));
 sg13g2_and2_1 _11241_ (.A(net1161),
    .B(_00925_),
    .X(_05247_));
 sg13g2_a22oi_1 _11242_ (.Y(_05248_),
    .B1(net1006),
    .B2(_05247_),
    .A2(_00923_),
    .A1(net958));
 sg13g2_and2_1 _11243_ (.A(net1161),
    .B(_00921_),
    .X(_05249_));
 sg13g2_a22oi_1 _11244_ (.Y(_05250_),
    .B1(net1004),
    .B2(_05249_),
    .A2(_00919_),
    .A1(net958));
 sg13g2_and2_1 _11245_ (.A(net1162),
    .B(_00924_),
    .X(_05251_));
 sg13g2_a22oi_1 _11246_ (.Y(_05252_),
    .B1(net1009),
    .B2(_05251_),
    .A2(_00922_),
    .A1(net958));
 sg13g2_nor4_1 _11247_ (.A(net916),
    .B(_05248_),
    .C(_05250_),
    .D(_05252_),
    .Y(_05253_));
 sg13g2_o21ai_1 _11248_ (.B1(_05253_),
    .Y(_05254_),
    .A1(net1001),
    .A2(_05246_));
 sg13g2_mux4_1 _11249_ (.S0(net1162),
    .A0(_00911_),
    .A1(_00913_),
    .A2(_00915_),
    .A3(_00917_),
    .S1(net1111),
    .X(_05255_));
 sg13g2_nand2_1 _11250_ (.Y(_05256_),
    .A(net1214),
    .B(_05255_));
 sg13g2_mux4_1 _11251_ (.S0(net1146),
    .A0(_00910_),
    .A1(_00912_),
    .A2(_00914_),
    .A3(_00916_),
    .S1(net1108),
    .X(_05257_));
 sg13g2_nand2_1 _11252_ (.Y(_05258_),
    .A(net972),
    .B(_05257_));
 sg13g2_a22oi_1 _11253_ (.Y(_05259_),
    .B1(net1402),
    .B2(net946),
    .A2(_05258_),
    .A1(_05256_));
 sg13g2_mux4_1 _11254_ (.S0(net1146),
    .A0(_00898_),
    .A1(_00900_),
    .A2(_00899_),
    .A3(_00901_),
    .S1(net1214),
    .X(_05260_));
 sg13g2_and2_1 _11255_ (.A(_04472_),
    .B(_05260_),
    .X(_05261_));
 sg13g2_nand2_1 _11256_ (.Y(_05262_),
    .A(net1173),
    .B(_00896_));
 sg13g2_nor2b_1 _11257_ (.A(net1176),
    .B_N(_00895_),
    .Y(_05263_));
 sg13g2_a22oi_1 _11258_ (.Y(_05264_),
    .B1(_05263_),
    .B2(net977),
    .A2(_00897_),
    .A1(net1176));
 sg13g2_a22oi_1 _11259_ (.Y(_05265_),
    .B1(_05264_),
    .B2(_04823_),
    .A2(_05262_),
    .A1(net976));
 sg13g2_nor4_1 _11260_ (.A(net895),
    .B(_05259_),
    .C(_05261_),
    .D(_05265_),
    .Y(_05266_));
 sg13g2_nor2_1 _11261_ (.A(net960),
    .B(_00904_),
    .Y(_05267_));
 sg13g2_nor2_1 _11262_ (.A(net1172),
    .B(_00902_),
    .Y(_05268_));
 sg13g2_a21oi_1 _11263_ (.A1(net935),
    .A2(_05267_),
    .Y(_05269_),
    .B1(_05268_));
 sg13g2_nor2b_1 _11264_ (.A(net1147),
    .B_N(_00906_),
    .Y(_05270_));
 sg13g2_a22oi_1 _11265_ (.Y(_05271_),
    .B1(net1009),
    .B2(_05270_),
    .A2(_00908_),
    .A1(net1172));
 sg13g2_mux4_1 _11266_ (.S0(net1172),
    .A0(_00903_),
    .A1(_00905_),
    .A2(_00907_),
    .A3(_00909_),
    .S1(net1108),
    .X(_05272_));
 sg13g2_nor2_1 _11267_ (.A(net973),
    .B(_05272_),
    .Y(_05273_));
 sg13g2_a22oi_1 _11268_ (.Y(_05274_),
    .B1(_05273_),
    .B2(net947),
    .A2(_05271_),
    .A1(net928));
 sg13g2_o21ai_1 _11269_ (.B1(_05274_),
    .Y(_05275_),
    .A1(net1000),
    .A2(_05269_));
 sg13g2_and3_1 _11270_ (.X(_05276_),
    .A(_05254_),
    .B(_05266_),
    .C(_05275_));
 sg13g2_buf_2 fanout660 (.A(net662),
    .X(net660));
 sg13g2_buf_1 fanout659 (.A(_02444_),
    .X(net659));
 sg13g2_and2_1 _11273_ (.A(_03547_),
    .B(net911),
    .X(_05279_));
 sg13g2_nand3_1 _11274_ (.B(_02572_),
    .C(net940),
    .A(net1260),
    .Y(_05280_));
 sg13g2_buf_2 fanout658 (.A(net659),
    .X(net658));
 sg13g2_a21oi_1 _11276_ (.A1(net3),
    .A2(net99),
    .Y(_05282_),
    .B1(_03837_));
 sg13g2_and3_1 _11277_ (.X(_05283_),
    .A(net901),
    .B(_05280_),
    .C(_05282_));
 sg13g2_or2_1 _11278_ (.X(_05284_),
    .B(_03836_),
    .A(net1261));
 sg13g2_inv_1 _11279_ (.Y(_05285_),
    .A(net1247));
 sg13g2_nand2_1 _11280_ (.Y(_05286_),
    .A(_05285_),
    .B(_02570_));
 sg13g2_a22oi_1 _11281_ (.Y(_05287_),
    .B1(net985),
    .B2(_03814_),
    .A2(_05286_),
    .A1(_05284_));
 sg13g2_a22oi_1 _11282_ (.Y(_05288_),
    .B1(_05283_),
    .B2(_05287_),
    .A2(_05279_),
    .A1(_03574_));
 sg13g2_buf_2 fanout657 (.A(net658),
    .X(net657));
 sg13g2_xnor2_1 _11284_ (.Y(_05290_),
    .A(net876),
    .B(net609));
 sg13g2_and2_1 _11285_ (.A(net611),
    .B(_05290_),
    .X(_05291_));
 sg13g2_buf_2 fanout656 (.A(net657),
    .X(net656));
 sg13g2_mux4_1 _11287_ (.S0(net1186),
    .A0(_00866_),
    .A1(_00868_),
    .A2(_00867_),
    .A3(_00869_),
    .S1(net1230),
    .X(_05293_));
 sg13g2_nor2_1 _11288_ (.A(net961),
    .B(_05293_),
    .Y(_05294_));
 sg13g2_mux2_1 _11289_ (.A0(_00863_),
    .A1(_00865_),
    .S(net1183),
    .X(_05295_));
 sg13g2_o21ai_1 _11290_ (.B1(_04577_),
    .Y(_05296_),
    .A1(net1005),
    .A2(_05295_));
 sg13g2_o21ai_1 _11291_ (.B1(net937),
    .Y(_05297_),
    .A1(_05294_),
    .A2(_05296_));
 sg13g2_nand2b_1 _11292_ (.Y(_05298_),
    .B(_03783_),
    .A_N(_00862_));
 sg13g2_or3_1 _11293_ (.A(_00864_),
    .B(net921),
    .C(_03790_),
    .X(_05299_));
 sg13g2_nand3_1 _11294_ (.B(_05298_),
    .C(_05299_),
    .A(_05297_),
    .Y(_05300_));
 sg13g2_mux4_1 _11295_ (.S0(net1186),
    .A0(_00890_),
    .A1(_00892_),
    .A2(_00891_),
    .A3(_00893_),
    .S1(net1230),
    .X(_05301_));
 sg13g2_mux4_1 _11296_ (.S0(net1181),
    .A0(_00886_),
    .A1(_00888_),
    .A2(_00887_),
    .A3(_00889_),
    .S1(net1230),
    .X(_05302_));
 sg13g2_mux2_1 _11297_ (.A0(_05301_),
    .A1(_05302_),
    .S(net961),
    .X(_05303_));
 sg13g2_mux4_1 _11298_ (.S0(net1186),
    .A0(_00879_),
    .A1(_00881_),
    .A2(_00883_),
    .A3(_00885_),
    .S1(net1116),
    .X(_05304_));
 sg13g2_mux4_1 _11299_ (.S0(net1186),
    .A0(_00878_),
    .A1(_00880_),
    .A2(_00882_),
    .A3(_00884_),
    .S1(net1116),
    .X(_05305_));
 sg13g2_mux2_1 _11300_ (.A0(_05304_),
    .A1(_05305_),
    .S(net981),
    .X(_05306_));
 sg13g2_a221oi_1 _11301_ (.B2(_04791_),
    .C1(net895),
    .B1(_05306_),
    .A1(net993),
    .Y(_05307_),
    .A2(_05303_));
 sg13g2_nor2b_1 _11302_ (.A(net1183),
    .B_N(_00874_),
    .Y(_05308_));
 sg13g2_a22oi_1 _11303_ (.Y(_05309_),
    .B1(_04518_),
    .B2(_05308_),
    .A2(_00876_),
    .A1(net1183));
 sg13g2_nor3_1 _11304_ (.A(net959),
    .B(_00872_),
    .C(net998),
    .Y(_05310_));
 sg13g2_mux4_1 _11305_ (.S0(net1186),
    .A0(_00871_),
    .A1(_00873_),
    .A2(_00875_),
    .A3(_00877_),
    .S1(net1114),
    .X(_05311_));
 sg13g2_nor2_1 _11306_ (.A(net977),
    .B(_05311_),
    .Y(_05312_));
 sg13g2_nor3_1 _11307_ (.A(net1183),
    .B(_00870_),
    .C(net998),
    .Y(_05313_));
 sg13g2_a22oi_1 _11308_ (.Y(_05314_),
    .B1(_05312_),
    .B2(_05313_),
    .A2(_05310_),
    .A1(net937));
 sg13g2_nand3b_1 _11309_ (.B(_05314_),
    .C(_04804_),
    .Y(_05315_),
    .A_N(_05309_));
 sg13g2_nand3_1 _11310_ (.B(_05307_),
    .C(_05315_),
    .A(_05300_),
    .Y(_05316_));
 sg13g2_buf_2 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_1 fanout654 (.A(net659),
    .X(net654));
 sg13g2_nand2_1 _11313_ (.Y(_05319_),
    .A(net18),
    .B(net943));
 sg13g2_nor2_1 _11314_ (.A(net909),
    .B(_05319_),
    .Y(_05320_));
 sg13g2_a21oi_1 _11315_ (.A1(net160),
    .A2(net908),
    .Y(_05321_),
    .B1(_05320_));
 sg13g2_xnor2_1 _11316_ (.Y(_05322_),
    .A(net874),
    .B(_05321_));
 sg13g2_buf_1 fanout653 (.A(net654),
    .X(net653));
 sg13g2_nor2_1 _11318_ (.A(net604),
    .B(_05322_),
    .Y(_05324_));
 sg13g2_nand2_1 _11319_ (.Y(_05325_),
    .A(net604),
    .B(_05322_));
 sg13g2_o21ai_1 _11320_ (.B1(_05325_),
    .Y(_05326_),
    .A1(_05291_),
    .A2(_05324_));
 sg13g2_a21oi_1 _11321_ (.A1(_03621_),
    .A2(_03650_),
    .Y(_05327_),
    .B1(net902));
 sg13g2_nand2_1 _11322_ (.Y(_05328_),
    .A(net20),
    .B(net933));
 sg13g2_nor2_1 _11323_ (.A(net910),
    .B(_05328_),
    .Y(_05329_));
 sg13g2_o21ai_1 _11324_ (.B1(net881),
    .Y(_05330_),
    .A1(_05327_),
    .A2(_05329_));
 sg13g2_or3_1 _11325_ (.A(net881),
    .B(_05327_),
    .C(_05329_),
    .X(_05331_));
 sg13g2_buf_2 fanout652 (.A(net653),
    .X(net652));
 sg13g2_and2_1 _11327_ (.A(_05330_),
    .B(_05331_),
    .X(_05333_));
 sg13g2_buf_2 fanout651 (.A(net654),
    .X(net651));
 sg13g2_nor2_1 _11329_ (.A(net960),
    .B(_00824_),
    .Y(_05335_));
 sg13g2_nor2_1 _11330_ (.A(net1187),
    .B(_00822_),
    .Y(_05336_));
 sg13g2_a21oi_1 _11331_ (.A1(net937),
    .A2(_05335_),
    .Y(_05337_),
    .B1(_05336_));
 sg13g2_mux4_1 _11332_ (.S0(net1182),
    .A0(_00826_),
    .A1(_00828_),
    .A2(_00827_),
    .A3(_00829_),
    .S1(net1229),
    .X(_05338_));
 sg13g2_inv_1 _11333_ (.Y(_05339_),
    .A(_05338_));
 sg13g2_and2_1 _11334_ (.A(net1182),
    .B(_00825_),
    .X(_05340_));
 sg13g2_a22oi_1 _11335_ (.Y(_05341_),
    .B1(net1005),
    .B2(_05340_),
    .A2(_00823_),
    .A1(net960));
 sg13g2_a22oi_1 _11336_ (.Y(_05342_),
    .B1(_05341_),
    .B2(net916),
    .A2(_05339_),
    .A1(net1116));
 sg13g2_o21ai_1 _11337_ (.B1(_05342_),
    .Y(_05343_),
    .A1(net999),
    .A2(_05337_));
 sg13g2_mux4_1 _11338_ (.S0(net1187),
    .A0(_00814_),
    .A1(_00816_),
    .A2(_00815_),
    .A3(_00817_),
    .S1(net1229),
    .X(_05344_));
 sg13g2_mux4_1 _11339_ (.S0(net1182),
    .A0(_00818_),
    .A1(_00820_),
    .A2(_00819_),
    .A3(_00821_),
    .S1(net1229),
    .X(_05345_));
 sg13g2_a221oi_1 _11340_ (.B2(net925),
    .C1(net895),
    .B1(_05345_),
    .A1(net914),
    .Y(_05346_),
    .A2(_05344_));
 sg13g2_mux4_1 _11341_ (.S0(net1176),
    .A0(_00810_),
    .A1(_00812_),
    .A2(_00811_),
    .A3(_00813_),
    .S1(net1226),
    .X(_05347_));
 sg13g2_nor2b_1 _11342_ (.A(_04014_),
    .B_N(_05347_),
    .Y(_05348_));
 sg13g2_o21ai_1 _11343_ (.B1(_00798_),
    .Y(_05349_),
    .A1(net977),
    .A2(_00799_));
 sg13g2_nor3_1 _11344_ (.A(net1400),
    .B(_04410_),
    .C(_05349_),
    .Y(_05350_));
 sg13g2_o21ai_1 _11345_ (.B1(net996),
    .Y(_05351_),
    .A1(_05348_),
    .A2(_05350_));
 sg13g2_mux4_1 _11346_ (.S0(net1175),
    .A0(_00802_),
    .A1(_00804_),
    .A2(_00803_),
    .A3(_00805_),
    .S1(net1226),
    .X(_05352_));
 sg13g2_nor2b_1 _11347_ (.A(net1400),
    .B_N(_00799_),
    .Y(_05353_));
 sg13g2_a22oi_1 _11348_ (.Y(_05354_),
    .B1(net990),
    .B2(_05353_),
    .A2(_00807_),
    .A1(net1400));
 sg13g2_mux2_1 _11349_ (.A0(_00801_),
    .A1(_00809_),
    .S(net1399),
    .X(_05355_));
 sg13g2_o21ai_1 _11350_ (.B1(_04312_),
    .Y(_05356_),
    .A1(net987),
    .A2(_05355_));
 sg13g2_mux2_1 _11351_ (.A0(_00800_),
    .A1(_00808_),
    .S(net1400),
    .X(_05357_));
 sg13g2_nor2b_1 _11352_ (.A(net1175),
    .B_N(net1400),
    .Y(_05358_));
 sg13g2_a221oi_1 _11353_ (.B2(_00806_),
    .C1(net1231),
    .B1(_05358_),
    .A1(net1175),
    .Y(_05359_),
    .A2(_05357_));
 sg13g2_nor4_1 _11354_ (.A(net921),
    .B(_05354_),
    .C(_05356_),
    .D(_05359_),
    .Y(_05360_));
 sg13g2_a21oi_1 _11355_ (.A1(_05123_),
    .A2(_05352_),
    .Y(_05361_),
    .B1(_05360_));
 sg13g2_and4_2 _11356_ (.A(_05343_),
    .B(_05346_),
    .C(_05351_),
    .D(_05361_),
    .X(_05362_));
 sg13g2_buf_1 fanout650 (.A(net654),
    .X(net650));
 sg13g2_nor2_1 _11358_ (.A(_04168_),
    .B(net923),
    .Y(_05364_));
 sg13g2_nor2_1 _11359_ (.A(net910),
    .B(_05364_),
    .Y(_05365_));
 sg13g2_a22oi_1 _11360_ (.Y(_05366_),
    .B1(_05365_),
    .B2(net877),
    .A2(net910),
    .A1(_03613_));
 sg13g2_buf_2 fanout649 (.A(net654),
    .X(net649));
 sg13g2_nand2_1 _11362_ (.Y(_05368_),
    .A(net19),
    .B(net940));
 sg13g2_nor2_1 _11363_ (.A(net910),
    .B(_05368_),
    .Y(_05369_));
 sg13g2_a22oi_1 _11364_ (.Y(_05370_),
    .B1(_05369_),
    .B2(net881),
    .A2(net910),
    .A1(net161));
 sg13g2_buf_2 fanout648 (.A(_03794_),
    .X(net648));
 sg13g2_nor2_1 _11366_ (.A(net959),
    .B(_00856_),
    .Y(_05372_));
 sg13g2_nor2_1 _11367_ (.A(net1181),
    .B(_00854_),
    .Y(_05373_));
 sg13g2_a22oi_1 _11368_ (.Y(_05374_),
    .B1(_05373_),
    .B2(net1115),
    .A2(_05372_),
    .A1(net937));
 sg13g2_and2_1 _11369_ (.A(net1181),
    .B(_00860_),
    .X(_05375_));
 sg13g2_a21oi_1 _11370_ (.A1(net959),
    .A2(_00858_),
    .Y(_05376_),
    .B1(_05375_));
 sg13g2_o21ai_1 _11371_ (.B1(net981),
    .Y(_05377_),
    .A1(net962),
    .A2(_05376_));
 sg13g2_mux4_1 _11372_ (.S0(net1181),
    .A0(_00855_),
    .A1(_00857_),
    .A2(_00859_),
    .A3(_00861_),
    .S1(net1115),
    .X(_05378_));
 sg13g2_inv_1 _11373_ (.Y(_05379_),
    .A(_05378_));
 sg13g2_a21oi_1 _11374_ (.A1(net1228),
    .A2(_05379_),
    .Y(_05380_),
    .B1(net916));
 sg13g2_o21ai_1 _11375_ (.B1(_05380_),
    .Y(_05381_),
    .A1(_05374_),
    .A2(_05377_));
 sg13g2_inv_1 _11376_ (.Y(_05382_),
    .A(_00848_));
 sg13g2_o21ai_1 _11377_ (.B1(_05382_),
    .Y(_05383_),
    .A1(net1034),
    .A2(net1020));
 sg13g2_mux4_1 _11378_ (.S0(net977),
    .A0(_00847_),
    .A1(_00846_),
    .A2(_00849_),
    .A3(_05383_),
    .S1(net1181),
    .X(_05384_));
 sg13g2_nand3_1 _11379_ (.B(net914),
    .C(_05384_),
    .A(net937),
    .Y(_05385_));
 sg13g2_and2_1 _11380_ (.A(net937),
    .B(net925),
    .X(_05386_));
 sg13g2_buf_2 fanout647 (.A(net648),
    .X(net647));
 sg13g2_inv_1 _11382_ (.Y(_05388_),
    .A(_00852_));
 sg13g2_o21ai_1 _11383_ (.B1(_05388_),
    .Y(_05389_),
    .A1(net1034),
    .A2(net1020));
 sg13g2_mux4_1 _11384_ (.S0(net977),
    .A0(_00851_),
    .A1(_00850_),
    .A2(_00853_),
    .A3(_05389_),
    .S1(net1181),
    .X(_05390_));
 sg13g2_nand2_1 _11385_ (.Y(_05391_),
    .A(_05386_),
    .B(_05390_));
 sg13g2_nor2b_1 _11386_ (.A(net1179),
    .B_N(_00842_),
    .Y(_05392_));
 sg13g2_a22oi_1 _11387_ (.Y(_05393_),
    .B1(net1008),
    .B2(_05392_),
    .A2(_00844_),
    .A1(net1179));
 sg13g2_mux4_1 _11388_ (.S0(net1178),
    .A0(_00839_),
    .A1(_00841_),
    .A2(_00843_),
    .A3(_00845_),
    .S1(net1114),
    .X(_05394_));
 sg13g2_nor2_1 _11389_ (.A(net977),
    .B(_05394_),
    .Y(_05395_));
 sg13g2_nor3_1 _11390_ (.A(net947),
    .B(_05393_),
    .C(_05395_),
    .Y(_05396_));
 sg13g2_or2_1 _11391_ (.X(_05397_),
    .B(_00838_),
    .A(net1180));
 sg13g2_nor2b_1 _11392_ (.A(_00840_),
    .B_N(net1180),
    .Y(_05398_));
 sg13g2_o21ai_1 _11393_ (.B1(_05398_),
    .Y(_05399_),
    .A1(net1034),
    .A2(net1020));
 sg13g2_a21o_1 _11394_ (.A2(_05399_),
    .A1(_05397_),
    .B1(net998),
    .X(_05400_));
 sg13g2_mux4_1 _11395_ (.S0(net1179),
    .A0(_00834_),
    .A1(_00836_),
    .A2(_00835_),
    .A3(_00837_),
    .S1(net1227),
    .X(_05401_));
 sg13g2_and3_1 _11396_ (.X(_05402_),
    .A(net995),
    .B(net968),
    .C(_05401_));
 sg13g2_nand2_1 _11397_ (.Y(_05403_),
    .A(_00831_),
    .B(_00830_));
 sg13g2_a22oi_1 _11398_ (.Y(_05404_),
    .B1(_04410_),
    .B2(net988),
    .A2(_05403_),
    .A1(net1228));
 sg13g2_or3_1 _11399_ (.A(net921),
    .B(_05402_),
    .C(_05404_),
    .X(_05405_));
 sg13g2_mux2_1 _11400_ (.A0(_00831_),
    .A1(_00833_),
    .S(net1180),
    .X(_05406_));
 sg13g2_nand2_1 _11401_ (.Y(_05407_),
    .A(net1228),
    .B(_05406_));
 sg13g2_nand2_1 _11402_ (.Y(_05408_),
    .A(_00832_),
    .B(_04238_));
 sg13g2_a21oi_1 _11403_ (.A1(_05407_),
    .A2(_05408_),
    .Y(_05409_),
    .B1(_04823_));
 sg13g2_a22oi_1 _11404_ (.Y(_05410_),
    .B1(_05405_),
    .B2(_05409_),
    .A2(_05400_),
    .A1(_05396_));
 sg13g2_nand4_1 _11405_ (.B(_05385_),
    .C(_05391_),
    .A(_05381_),
    .Y(_05411_),
    .D(_05410_));
 sg13g2_buf_1 fanout646 (.A(_03843_),
    .X(net646));
 sg13g2_nor3_1 _11407_ (.A(_05366_),
    .B(_05370_),
    .C(net602),
    .Y(_05413_));
 sg13g2_a21oi_1 _11408_ (.A1(_05333_),
    .A2(_05362_),
    .Y(_05414_),
    .B1(_05413_));
 sg13g2_o21ai_1 _11409_ (.B1(_05411_),
    .Y(_05415_),
    .A1(_05366_),
    .A2(_05370_));
 sg13g2_a21o_1 _11410_ (.A2(_05331_),
    .A1(_05330_),
    .B1(_05415_),
    .X(_05416_));
 sg13g2_and3_1 _11411_ (.X(_05417_),
    .A(_05330_),
    .B(_05331_),
    .C(_05415_));
 sg13g2_a21oi_1 _11412_ (.A1(_05362_),
    .A2(_05416_),
    .Y(_05418_),
    .B1(_05417_));
 sg13g2_a21o_1 _11413_ (.A2(_05414_),
    .A1(_05326_),
    .B1(_05418_),
    .X(_05419_));
 sg13g2_nand4_1 _11414_ (.B(_05346_),
    .C(_05351_),
    .A(_05343_),
    .Y(_05420_),
    .D(_05361_));
 sg13g2_buf_1 fanout645 (.A(net646),
    .X(net645));
 sg13g2_buf_2 fanout644 (.A(net645),
    .X(net644));
 sg13g2_xnor2_1 _11417_ (.Y(_05423_),
    .A(_05333_),
    .B(net601));
 sg13g2_buf_4 fanout643 (.X(net643),
    .A(net645));
 sg13g2_xnor2_1 _11419_ (.Y(_05425_),
    .A(net604),
    .B(_05322_));
 sg13g2_nor2_1 _11420_ (.A(_05366_),
    .B(_05370_),
    .Y(_05426_));
 sg13g2_and4_1 _11421_ (.A(_05381_),
    .B(_05385_),
    .C(_05391_),
    .D(_05410_),
    .X(_05427_));
 sg13g2_buf_4 fanout642 (.X(net642),
    .A(_03843_));
 sg13g2_xnor2_1 _11423_ (.Y(_05429_),
    .A(_05426_),
    .B(_05427_));
 sg13g2_nor2_1 _11424_ (.A(_05425_),
    .B(_05429_),
    .Y(_05430_));
 sg13g2_nand2_1 _11425_ (.Y(_05431_),
    .A(_05423_),
    .B(_05430_));
 sg13g2_nand2_1 _11426_ (.Y(_05432_),
    .A(_05419_),
    .B(_05431_));
 sg13g2_a21oi_1 _11427_ (.A1(_05326_),
    .A2(_05414_),
    .Y(_05433_),
    .B1(_05418_));
 sg13g2_nand3_1 _11428_ (.B(_05266_),
    .C(_05275_),
    .A(_05254_),
    .Y(_05434_));
 sg13g2_buf_1 fanout641 (.A(net642),
    .X(net641));
 sg13g2_xnor2_1 _11430_ (.Y(_05436_),
    .A(_05434_),
    .B(_05290_));
 sg13g2_o21ai_1 _11431_ (.B1(net909),
    .Y(_05437_),
    .A1(_03524_),
    .A2(_03541_));
 sg13g2_buf_1 fanout640 (.A(net641),
    .X(net640));
 sg13g2_nand3b_1 _11433_ (.B(net1251),
    .C(net1254),
    .Y(_05439_),
    .A_N(net1273));
 sg13g2_or3_1 _11434_ (.A(net1251),
    .B(net1254),
    .C(net1257),
    .X(_05440_));
 sg13g2_a22oi_1 _11435_ (.Y(_05441_),
    .B1(net985),
    .B2(_03814_),
    .A2(_05440_),
    .A1(_05439_));
 sg13g2_buf_2 fanout639 (.A(net640),
    .X(net639));
 sg13g2_nor2_1 _11437_ (.A(net1248),
    .B(net1257),
    .Y(_05443_));
 sg13g2_nand3_1 _11438_ (.B(net1254),
    .C(net1248),
    .A(net1251),
    .Y(_05444_));
 sg13g2_o21ai_1 _11439_ (.B1(_05444_),
    .Y(_05445_),
    .A1(net986),
    .A2(_05443_));
 sg13g2_nor2_1 _11440_ (.A(_03812_),
    .B(_03829_),
    .Y(_05446_));
 sg13g2_nand3b_1 _11441_ (.B(_05445_),
    .C(_05446_),
    .Y(_05447_),
    .A_N(_05441_));
 sg13g2_xnor2_1 _11442_ (.Y(_05448_),
    .A(net1252),
    .B(net1255));
 sg13g2_nand3_1 _11443_ (.B(_03824_),
    .C(_05448_),
    .A(_02561_),
    .Y(_05449_));
 sg13g2_buf_1 fanout638 (.A(_03877_),
    .X(net638));
 sg13g2_nand3_1 _11445_ (.B(net940),
    .C(_05449_),
    .A(_02572_),
    .Y(_05451_));
 sg13g2_a21oi_1 _11446_ (.A1(_05446_),
    .A2(_05445_),
    .Y(_05452_),
    .B1(net1273));
 sg13g2_a221oi_1 _11447_ (.B2(_05451_),
    .C1(_05452_),
    .B1(_05447_),
    .A1(_03127_),
    .Y(_05453_),
    .A2(_05441_));
 sg13g2_buf_1 fanout637 (.A(net638),
    .X(net637));
 sg13g2_nand2_2 _11449_ (.Y(_05455_),
    .A(net902),
    .B(net871));
 sg13g2_nand2_1 _11450_ (.Y(_05456_),
    .A(_05437_),
    .B(_05455_));
 sg13g2_buf_2 fanout636 (.A(net638),
    .X(net636));
 sg13g2_xnor2_1 _11452_ (.Y(_05458_),
    .A(net874),
    .B(net400));
 sg13g2_mux4_1 _11453_ (.S0(net1200),
    .A0(_00946_),
    .A1(_00948_),
    .A2(_00947_),
    .A3(_00949_),
    .S1(net1232),
    .X(_05459_));
 sg13g2_nand3_1 _11454_ (.B(_03749_),
    .C(_05061_),
    .A(_00954_),
    .Y(_05460_));
 sg13g2_a21oi_1 _11455_ (.A1(net1198),
    .A2(_00956_),
    .Y(_05461_),
    .B1(net1232));
 sg13g2_or2_1 _11456_ (.X(_05462_),
    .B(_05461_),
    .A(_05064_));
 sg13g2_nor2b_1 _11457_ (.A(net1198),
    .B_N(_00955_),
    .Y(_05463_));
 sg13g2_a22oi_1 _11458_ (.Y(_05464_),
    .B1(_05463_),
    .B2(net979),
    .A2(_00957_),
    .A1(net1198));
 sg13g2_a22oi_1 _11459_ (.Y(_05465_),
    .B1(_05464_),
    .B2(net922),
    .A2(_05462_),
    .A1(_05460_));
 sg13g2_a21oi_1 _11460_ (.A1(_05386_),
    .A2(_05459_),
    .Y(_05466_),
    .B1(_05465_));
 sg13g2_mux4_1 _11461_ (.S0(net1200),
    .A0(_00942_),
    .A1(_00944_),
    .A2(_00943_),
    .A3(_00945_),
    .S1(net1232),
    .X(_05467_));
 sg13g2_and2_1 _11462_ (.A(net914),
    .B(_05467_),
    .X(_05468_));
 sg13g2_nand3_1 _11463_ (.B(net993),
    .C(_05073_),
    .A(_00950_),
    .Y(_05469_));
 sg13g2_a21oi_1 _11464_ (.A1(net1199),
    .A2(_00952_),
    .Y(_05470_),
    .B1(net1232));
 sg13g2_or2_1 _11465_ (.X(_05471_),
    .B(_05470_),
    .A(_05075_));
 sg13g2_nor2b_1 _11466_ (.A(net1199),
    .B_N(_00951_),
    .Y(_05472_));
 sg13g2_a22oi_1 _11467_ (.Y(_05473_),
    .B1(_05472_),
    .B2(net979),
    .A2(_00953_),
    .A1(net1199));
 sg13g2_a21oi_1 _11468_ (.A1(_05469_),
    .A2(_05471_),
    .Y(_05474_),
    .B1(_05473_));
 sg13g2_o21ai_1 _11469_ (.B1(net943),
    .Y(_05475_),
    .A1(_05468_),
    .A2(_05474_));
 sg13g2_nor2b_1 _11470_ (.A(net1198),
    .B_N(_00930_),
    .Y(_05476_));
 sg13g2_a22oi_1 _11471_ (.Y(_05477_),
    .B1(net1010),
    .B2(_05476_),
    .A2(_00932_),
    .A1(net1199));
 sg13g2_nor2b_1 _11472_ (.A(net1120),
    .B_N(_00927_),
    .Y(_05478_));
 sg13g2_a22oi_1 _11473_ (.Y(_05479_),
    .B1(net990),
    .B2(_05478_),
    .A2(_00931_),
    .A1(net1120));
 sg13g2_nor2b_1 _11474_ (.A(net1120),
    .B_N(_00929_),
    .Y(_05480_));
 sg13g2_a22oi_1 _11475_ (.Y(_05481_),
    .B1(net987),
    .B2(_05480_),
    .A2(_00933_),
    .A1(net1120));
 sg13g2_nand2b_1 _11476_ (.Y(_05482_),
    .B(net1201),
    .A_N(_00928_));
 sg13g2_o21ai_1 _11477_ (.B1(_04577_),
    .Y(_05483_),
    .A1(net1000),
    .A2(_05482_));
 sg13g2_nor4_1 _11478_ (.A(_05477_),
    .B(_05479_),
    .C(_05481_),
    .D(_05483_),
    .Y(_05484_));
 sg13g2_nand2b_1 _11479_ (.Y(_05485_),
    .B(_03783_),
    .A_N(_00926_));
 sg13g2_o21ai_1 _11480_ (.B1(_05485_),
    .Y(_05486_),
    .A1(net923),
    .A2(_05484_));
 sg13g2_or3_1 _11481_ (.A(_00936_),
    .B(net923),
    .C(_03790_),
    .X(_05487_));
 sg13g2_mux4_1 _11482_ (.S0(net1201),
    .A0(_00935_),
    .A1(_00937_),
    .A2(_00939_),
    .A3(_00941_),
    .S1(net1120),
    .X(_05488_));
 sg13g2_nand2b_1 _11483_ (.Y(_05489_),
    .B(net1233),
    .A_N(_05488_));
 sg13g2_or3_1 _11484_ (.A(net1201),
    .B(_00934_),
    .C(net1000),
    .X(_05490_));
 sg13g2_nand2b_1 _11485_ (.Y(_05491_),
    .B(net1201),
    .A_N(_00940_));
 sg13g2_o21ai_1 _11486_ (.B1(_05491_),
    .Y(_05492_),
    .A1(net1201),
    .A2(_00938_));
 sg13g2_a22oi_1 _11487_ (.Y(_05493_),
    .B1(net922),
    .B2(_05137_),
    .A2(_05492_),
    .A1(_03935_));
 sg13g2_nand4_1 _11488_ (.B(_05489_),
    .C(_05490_),
    .A(_05487_),
    .Y(_05494_),
    .D(_05493_));
 sg13g2_and4_1 _11489_ (.A(_05466_),
    .B(_05475_),
    .C(_05486_),
    .D(_05494_),
    .X(_05495_));
 sg13g2_buf_2 fanout635 (.A(net638),
    .X(net635));
 sg13g2_buf_2 fanout634 (.A(net635),
    .X(net634));
 sg13g2_and2_1 _11492_ (.A(_03747_),
    .B(net597),
    .X(_05498_));
 sg13g2_buf_1 fanout633 (.A(_04101_),
    .X(net633));
 sg13g2_nand3_1 _11494_ (.B(_05458_),
    .C(_05498_),
    .A(_05436_),
    .Y(_05500_));
 sg13g2_buf_2 fanout632 (.A(_04101_),
    .X(net632));
 sg13g2_nor2_1 _11496_ (.A(net1248),
    .B(net32),
    .Y(_05502_));
 sg13g2_o21ai_1 _11497_ (.B1(_05444_),
    .Y(_05503_),
    .A1(net986),
    .A2(_05502_));
 sg13g2_nand2_1 _11498_ (.Y(_05504_),
    .A(_05446_),
    .B(_05503_));
 sg13g2_nand4_1 _11499_ (.B(_02572_),
    .C(net941),
    .A(net1277),
    .Y(_05505_),
    .D(_05449_));
 sg13g2_buf_2 fanout631 (.A(_04166_),
    .X(net631));
 sg13g2_nand2b_1 _11501_ (.Y(_05507_),
    .B(_03127_),
    .A_N(_03836_));
 sg13g2_inv_1 _11502_ (.Y(_05508_),
    .A(net1244));
 sg13g2_nand2_1 _11503_ (.Y(_05509_),
    .A(_05508_),
    .B(_02570_));
 sg13g2_a22oi_1 _11504_ (.Y(_05510_),
    .B1(net985),
    .B2(_03814_),
    .A2(_05509_),
    .A1(_05507_));
 sg13g2_a22oi_1 _11505_ (.Y(_05511_),
    .B1(net908),
    .B2(_05510_),
    .A2(_05505_),
    .A1(_05504_));
 sg13g2_a21o_1 _11506_ (.A2(net908),
    .A1(net155),
    .B1(_05511_),
    .X(_05512_));
 sg13g2_buf_1 fanout630 (.A(_04343_),
    .X(net630));
 sg13g2_buf_2 fanout629 (.A(_04343_),
    .X(net629));
 sg13g2_a22oi_1 _11509_ (.Y(_05515_),
    .B1(net390),
    .B2(net598),
    .A2(_05455_),
    .A1(_05437_));
 sg13g2_a21oi_1 _11510_ (.A1(net155),
    .A2(net908),
    .Y(_05516_),
    .B1(_05511_));
 sg13g2_buf_2 fanout628 (.A(net629),
    .X(net628));
 sg13g2_a21o_1 _11512_ (.A2(_03523_),
    .A1(_03514_),
    .B1(_03127_),
    .X(_05518_));
 sg13g2_nor2_1 _11513_ (.A(_03531_),
    .B(_03540_),
    .Y(_05519_));
 sg13g2_a21oi_2 _11514_ (.B1(net901),
    .Y(_05520_),
    .A2(_05519_),
    .A1(_05518_));
 sg13g2_and2_1 _11515_ (.A(net901),
    .B(net871),
    .X(_05521_));
 sg13g2_buf_2 fanout627 (.A(net628),
    .X(net627));
 sg13g2_nor4_1 _11517_ (.A(net377),
    .B(net598),
    .C(_05520_),
    .D(_05521_),
    .Y(_05523_));
 sg13g2_nor4_1 _11518_ (.A(net882),
    .B(net389),
    .C(_05520_),
    .D(_05521_),
    .Y(_05524_));
 sg13g2_a22oi_1 _11519_ (.Y(_05525_),
    .B1(net874),
    .B2(net377),
    .A2(_05455_),
    .A1(_05437_));
 sg13g2_nor4_1 _11520_ (.A(_05515_),
    .B(_05523_),
    .C(_05524_),
    .D(_05525_),
    .Y(_05526_));
 sg13g2_inv_1 _11521_ (.Y(_05527_),
    .A(_00962_));
 sg13g2_a22oi_1 _11522_ (.Y(_05528_),
    .B1(net988),
    .B2(net1234),
    .A2(_05061_),
    .A1(_05527_));
 sg13g2_nand2b_1 _11523_ (.Y(_05529_),
    .B(_00960_),
    .A_N(net1121));
 sg13g2_nand2_1 _11524_ (.Y(_05530_),
    .A(net1121),
    .B(_00964_));
 sg13g2_nand3_1 _11525_ (.B(_05529_),
    .C(_05530_),
    .A(net1198),
    .Y(_05531_));
 sg13g2_a21o_1 _11526_ (.A2(_05531_),
    .A1(_05528_),
    .B1(net923),
    .X(_05532_));
 sg13g2_a21o_1 _11527_ (.A2(_04410_),
    .A1(net942),
    .B1(_00958_),
    .X(_05533_));
 sg13g2_and2_1 _11528_ (.A(_05532_),
    .B(_05533_),
    .X(_05534_));
 sg13g2_buf_2 fanout626 (.A(_04389_),
    .X(net626));
 sg13g2_mux2_1 _11530_ (.A0(_00968_),
    .A1(_00972_),
    .S(net1117),
    .X(_05536_));
 sg13g2_nand2_1 _11531_ (.Y(_05537_),
    .A(_04238_),
    .B(_05536_));
 sg13g2_mux2_1 _11532_ (.A0(_00966_),
    .A1(_00970_),
    .S(net1117),
    .X(_05538_));
 sg13g2_nand2_1 _11533_ (.Y(_05539_),
    .A(_03743_),
    .B(_05538_));
 sg13g2_a21oi_1 _11534_ (.A1(_05537_),
    .A2(_05539_),
    .Y(_05540_),
    .B1(net948));
 sg13g2_mux4_1 _11535_ (.S0(net1200),
    .A0(_00978_),
    .A1(_00980_),
    .A2(_00979_),
    .A3(_00981_),
    .S1(net1233),
    .X(_05541_));
 sg13g2_nand3_1 _11536_ (.B(_03737_),
    .C(_05541_),
    .A(net943),
    .Y(_05542_));
 sg13g2_mux4_1 _11537_ (.S0(net1199),
    .A0(_00982_),
    .A1(_00984_),
    .A2(_00983_),
    .A3(_00985_),
    .S1(net1232),
    .X(_05543_));
 sg13g2_nand4_1 _11538_ (.B(net943),
    .C(_03756_),
    .A(net1394),
    .Y(_05544_),
    .D(_05543_));
 sg13g2_nand3b_1 _11539_ (.B(_05542_),
    .C(_05544_),
    .Y(_05545_),
    .A_N(_05540_));
 sg13g2_buf_2 fanout625 (.A(_04486_),
    .X(net625));
 sg13g2_mux2_1 _11541_ (.A0(_00965_),
    .A1(_00973_),
    .S(net1401),
    .X(_05547_));
 sg13g2_mux2_1 _11542_ (.A0(_00963_),
    .A1(_00971_),
    .S(net1401),
    .X(_05548_));
 sg13g2_mux2_1 _11543_ (.A0(_00961_),
    .A1(_00969_),
    .S(net1402),
    .X(_05549_));
 sg13g2_mux2_1 _11544_ (.A0(_00959_),
    .A1(_00967_),
    .S(net1402),
    .X(_05550_));
 sg13g2_mux4_1 _11545_ (.S0(net960),
    .A0(_05547_),
    .A1(_05548_),
    .A2(_05549_),
    .A3(_05550_),
    .S1(net962),
    .X(_05551_));
 sg13g2_and4_1 _11546_ (.A(net1233),
    .B(net997),
    .C(net942),
    .D(_05551_),
    .X(_05552_));
 sg13g2_mux4_1 _11547_ (.S0(net1202),
    .A0(_00974_),
    .A1(_00976_),
    .A2(_00975_),
    .A3(_00977_),
    .S1(net1233),
    .X(_05553_));
 sg13g2_and3_1 _11548_ (.X(_05554_),
    .A(net943),
    .B(net914),
    .C(_05553_));
 sg13g2_nand3_1 _11549_ (.B(net993),
    .C(_05061_),
    .A(_00986_),
    .Y(_05555_));
 sg13g2_a21oi_1 _11550_ (.A1(net1199),
    .A2(_00988_),
    .Y(_05556_),
    .B1(net1232));
 sg13g2_or2_1 _11551_ (.X(_05557_),
    .B(_05556_),
    .A(_05064_));
 sg13g2_nor2b_1 _11552_ (.A(net1198),
    .B_N(_00987_),
    .Y(_05558_));
 sg13g2_a22oi_1 _11553_ (.Y(_05559_),
    .B1(_05558_),
    .B2(net979),
    .A2(_00989_),
    .A1(net1198));
 sg13g2_a22oi_1 _11554_ (.Y(_05560_),
    .B1(_05559_),
    .B2(net922),
    .A2(_05557_),
    .A1(_05555_));
 sg13g2_or3_1 _11555_ (.A(_05552_),
    .B(_05554_),
    .C(_05560_),
    .X(_05561_));
 sg13g2_buf_2 fanout624 (.A(net625),
    .X(net624));
 sg13g2_nor4_2 _11557_ (.A(net895),
    .B(_05534_),
    .C(_05545_),
    .Y(_05563_),
    .D(_05561_));
 sg13g2_buf_2 fanout623 (.A(_04592_),
    .X(net623));
 sg13g2_nand3_1 _11559_ (.B(_05526_),
    .C(net596),
    .A(_05436_),
    .Y(_05565_));
 sg13g2_nand2_2 _11560_ (.Y(_05566_),
    .A(_05500_),
    .B(_05565_));
 sg13g2_a21oi_2 _11561_ (.B1(_05510_),
    .Y(_05567_),
    .A2(_05505_),
    .A1(_05504_));
 sg13g2_buf_1 fanout622 (.A(_04632_),
    .X(net622));
 sg13g2_nor2_1 _11563_ (.A(_05567_),
    .B(net871),
    .Y(_05569_));
 sg13g2_and2_1 _11564_ (.A(_05567_),
    .B(net871),
    .X(_05570_));
 sg13g2_nor3_1 _11565_ (.A(net155),
    .B(_03524_),
    .C(_03541_),
    .Y(_05571_));
 sg13g2_a21oi_1 _11566_ (.A1(_05518_),
    .A2(_05519_),
    .Y(_05572_),
    .B1(_03501_));
 sg13g2_mux4_1 _11567_ (.S0(net874),
    .A0(_05569_),
    .A1(_05570_),
    .A2(_05571_),
    .A3(_05572_),
    .S1(net908),
    .X(_05573_));
 sg13g2_nor2b_1 _11568_ (.A(net597),
    .B_N(_05573_),
    .Y(_05574_));
 sg13g2_nor2_1 _11569_ (.A(_05520_),
    .B(_05521_),
    .Y(_05575_));
 sg13g2_buf_2 fanout621 (.A(net622),
    .X(net621));
 sg13g2_and4_1 _11571_ (.A(net875),
    .B(net389),
    .C(net597),
    .D(net368),
    .X(_05577_));
 sg13g2_nand2_1 _11572_ (.Y(_05578_),
    .A(_05532_),
    .B(_05533_));
 sg13g2_nor2_1 _11573_ (.A(net922),
    .B(_05075_),
    .Y(_05579_));
 sg13g2_a221oi_1 _11574_ (.B2(_05543_),
    .C1(_05540_),
    .B1(_05579_),
    .A1(_05386_),
    .Y(_05580_),
    .A2(_05541_));
 sg13g2_buf_2 fanout620 (.A(_04780_),
    .X(net620));
 sg13g2_nor3_1 _11576_ (.A(_05552_),
    .B(_05554_),
    .C(_05560_),
    .Y(_05582_));
 sg13g2_nand3_1 _11577_ (.B(_05580_),
    .C(_05582_),
    .A(_05578_),
    .Y(_05583_));
 sg13g2_buf_1 fanout619 (.A(_04883_),
    .X(net619));
 sg13g2_o21ai_1 _11579_ (.B1(_05583_),
    .Y(_05585_),
    .A1(_05574_),
    .A2(_05577_));
 sg13g2_nand2_1 _11580_ (.Y(_05586_),
    .A(_04827_),
    .B(_05573_));
 sg13g2_a22oi_1 _11581_ (.Y(_05587_),
    .B1(net881),
    .B2(net389),
    .A2(_05455_),
    .A1(_05437_));
 sg13g2_nor4_1 _11582_ (.A(net875),
    .B(net377),
    .C(_05520_),
    .D(_05521_),
    .Y(_05588_));
 sg13g2_nor2_1 _11583_ (.A(net597),
    .B(_05583_),
    .Y(_05589_));
 sg13g2_o21ai_1 _11584_ (.B1(_05589_),
    .Y(_05590_),
    .A1(_05587_),
    .A2(_05588_));
 sg13g2_nor3_2 _11585_ (.A(_05534_),
    .B(_05545_),
    .C(_05561_),
    .Y(_05591_));
 sg13g2_nor2_1 _11586_ (.A(net874),
    .B(net377),
    .Y(_05592_));
 sg13g2_nand4_1 _11587_ (.B(net400),
    .C(_05591_),
    .A(net597),
    .Y(_05593_),
    .D(_05592_));
 sg13g2_a22oi_1 _11588_ (.Y(_05594_),
    .B1(_05591_),
    .B2(net875),
    .A2(_05455_),
    .A1(_05437_));
 sg13g2_nor4_1 _11589_ (.A(net881),
    .B(_05520_),
    .C(_05521_),
    .D(_05583_),
    .Y(_05595_));
 sg13g2_and2_1 _11590_ (.A(net377),
    .B(net597),
    .X(_05596_));
 sg13g2_o21ai_1 _11591_ (.B1(_05596_),
    .Y(_05597_),
    .A1(_05594_),
    .A2(_05595_));
 sg13g2_and4_1 _11592_ (.A(_05586_),
    .B(_05590_),
    .C(_05593_),
    .D(_05597_),
    .X(_05598_));
 sg13g2_a21o_2 _11593_ (.A2(net911),
    .A1(_03448_),
    .B1(_03842_),
    .X(_05599_));
 sg13g2_buf_2 fanout618 (.A(_04883_),
    .X(net618));
 sg13g2_nor2b_1 _11595_ (.A(net1117),
    .B_N(_00993_),
    .Y(_05601_));
 sg13g2_a22oi_1 _11596_ (.Y(_05602_),
    .B1(net987),
    .B2(_05601_),
    .A2(_00997_),
    .A1(net1118));
 sg13g2_nor2b_1 _11597_ (.A(net1194),
    .B_N(_00994_),
    .Y(_05603_));
 sg13g2_a22oi_1 _11598_ (.Y(_05604_),
    .B1(net1009),
    .B2(_05603_),
    .A2(_00996_),
    .A1(net1194));
 sg13g2_nor2b_1 _11599_ (.A(net1118),
    .B_N(_00991_),
    .Y(_05605_));
 sg13g2_a22oi_1 _11600_ (.Y(_05606_),
    .B1(net990),
    .B2(_05605_),
    .A2(_00995_),
    .A1(net1118));
 sg13g2_or4_1 _11601_ (.A(net988),
    .B(_05602_),
    .C(_05604_),
    .D(_05606_),
    .X(_05607_));
 sg13g2_nor3_1 _11602_ (.A(_00992_),
    .B(net922),
    .C(_03790_),
    .Y(_05608_));
 sg13g2_nor2b_1 _11603_ (.A(_00990_),
    .B_N(_03783_),
    .Y(_05609_));
 sg13g2_a22oi_1 _11604_ (.Y(_05610_),
    .B1(_05608_),
    .B2(_05609_),
    .A2(_05607_),
    .A1(net942));
 sg13g2_nor2b_1 _11605_ (.A(_01000_),
    .B_N(net1191),
    .Y(_05611_));
 sg13g2_o21ai_1 _11606_ (.B1(_05611_),
    .Y(_05612_),
    .A1(net1037),
    .A2(net1023));
 sg13g2_o21ai_1 _11607_ (.B1(_05612_),
    .Y(_05613_),
    .A1(net1192),
    .A2(_00998_));
 sg13g2_nor2b_1 _11608_ (.A(net1117),
    .B_N(_00999_),
    .Y(_05614_));
 sg13g2_a22oi_1 _11609_ (.Y(_05615_),
    .B1(net990),
    .B2(_05614_),
    .A2(_01003_),
    .A1(net1117));
 sg13g2_nor2b_1 _11610_ (.A(net1118),
    .B_N(_01001_),
    .Y(_05616_));
 sg13g2_a22oi_1 _11611_ (.Y(_05617_),
    .B1(net987),
    .B2(_05616_),
    .A2(_01005_),
    .A1(net1117));
 sg13g2_or3_1 _11612_ (.A(net948),
    .B(_05615_),
    .C(_05617_),
    .X(_05618_));
 sg13g2_nor2b_1 _11613_ (.A(net1192),
    .B_N(_01002_),
    .Y(_05619_));
 sg13g2_a22oi_1 _11614_ (.Y(_05620_),
    .B1(_04518_),
    .B2(_05619_),
    .A2(_01004_),
    .A1(net1192));
 sg13g2_a22oi_1 _11615_ (.Y(_05621_),
    .B1(_05618_),
    .B2(_05620_),
    .A2(_05613_),
    .A1(net1041));
 sg13g2_nand3_1 _11616_ (.B(net993),
    .C(_05073_),
    .A(_01014_),
    .Y(_05622_));
 sg13g2_a21oi_1 _11617_ (.A1(net1196),
    .A2(_01016_),
    .Y(_05623_),
    .B1(net1234));
 sg13g2_or2_1 _11618_ (.X(_05624_),
    .B(_05623_),
    .A(_05075_));
 sg13g2_nor2b_1 _11619_ (.A(net1196),
    .B_N(_01015_),
    .Y(_05625_));
 sg13g2_a22oi_1 _11620_ (.Y(_05626_),
    .B1(_05625_),
    .B2(net978),
    .A2(_01017_),
    .A1(net1197));
 sg13g2_a22oi_1 _11621_ (.Y(_05627_),
    .B1(_05626_),
    .B2(net922),
    .A2(_05624_),
    .A1(_05622_));
 sg13g2_nand3_1 _11622_ (.B(net993),
    .C(_05061_),
    .A(_01018_),
    .Y(_05628_));
 sg13g2_a21oi_1 _11623_ (.A1(net1196),
    .A2(_01020_),
    .Y(_05629_),
    .B1(net1234));
 sg13g2_or2_1 _11624_ (.X(_05630_),
    .B(_05629_),
    .A(_05064_));
 sg13g2_nor2b_1 _11625_ (.A(net1197),
    .B_N(_01019_),
    .Y(_05631_));
 sg13g2_a22oi_1 _11626_ (.Y(_05632_),
    .B1(_05631_),
    .B2(net978),
    .A2(_01021_),
    .A1(net1197));
 sg13g2_a22oi_1 _11627_ (.Y(_05633_),
    .B1(_05632_),
    .B2(net922),
    .A2(_05630_),
    .A1(_05628_));
 sg13g2_mux4_1 _11628_ (.S0(net1195),
    .A0(_01006_),
    .A1(_01008_),
    .A2(_01007_),
    .A3(_01009_),
    .S1(net1234),
    .X(_05634_));
 sg13g2_and3_1 _11629_ (.X(_05635_),
    .A(net942),
    .B(net915),
    .C(_05634_));
 sg13g2_mux4_1 _11630_ (.S0(net1196),
    .A0(_01010_),
    .A1(_01012_),
    .A2(_01011_),
    .A3(_01013_),
    .S1(net1234),
    .X(_05636_));
 sg13g2_and3_1 _11631_ (.X(_05637_),
    .A(net942),
    .B(_03737_),
    .C(_05636_));
 sg13g2_or4_1 _11632_ (.A(_05627_),
    .B(_05633_),
    .C(_05635_),
    .D(_05637_),
    .X(_05638_));
 sg13g2_or4_1 _11633_ (.A(_04827_),
    .B(_05610_),
    .C(_05621_),
    .D(_05638_),
    .X(_05639_));
 sg13g2_buf_2 fanout617 (.A(_04972_),
    .X(net617));
 sg13g2_nand3_1 _11635_ (.B(_02572_),
    .C(net940),
    .A(net1301),
    .Y(_05641_));
 sg13g2_buf_1 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_2 fanout615 (.A(net616),
    .X(net615));
 sg13g2_a21oi_1 _11638_ (.A1(net31),
    .A2(net99),
    .Y(_05644_),
    .B1(_03837_));
 sg13g2_inv_1 _11639_ (.Y(_05645_),
    .A(net31));
 sg13g2_nand3_1 _11640_ (.B(net1251),
    .C(net1254),
    .A(net1301),
    .Y(_05646_));
 sg13g2_o21ai_1 _11641_ (.B1(_05646_),
    .Y(_05647_),
    .A1(_05645_),
    .A2(net986));
 sg13g2_a21oi_1 _11642_ (.A1(_02565_),
    .A2(_05647_),
    .Y(_05648_),
    .B1(_05449_));
 sg13g2_a22oi_1 _11643_ (.Y(_05649_),
    .B1(_05648_),
    .B2(net908),
    .A2(_05644_),
    .A1(_05641_));
 sg13g2_a21oi_1 _11644_ (.A1(net144),
    .A2(net910),
    .Y(_05650_),
    .B1(_05649_));
 sg13g2_buf_1 fanout614 (.A(_05026_),
    .X(net614));
 sg13g2_nand2_1 _11646_ (.Y(_05652_),
    .A(net881),
    .B(net584));
 sg13g2_o21ai_1 _11647_ (.B1(_05652_),
    .Y(_05653_),
    .A1(net587),
    .A2(net584));
 sg13g2_a21o_1 _11648_ (.A2(net910),
    .A1(net144),
    .B1(_05649_),
    .X(_05654_));
 sg13g2_buf_2 fanout613 (.A(_05026_),
    .X(net613));
 sg13g2_nor3_2 _11650_ (.A(_05610_),
    .B(_05621_),
    .C(_05638_),
    .Y(_05656_));
 sg13g2_buf_2 fanout612 (.A(_05203_),
    .X(net612));
 sg13g2_a21oi_1 _11652_ (.A1(net874),
    .A2(net575),
    .Y(_05658_),
    .B1(_05656_));
 sg13g2_o21ai_1 _11653_ (.B1(_05652_),
    .Y(_05659_),
    .A1(net594),
    .A2(_05658_));
 sg13g2_xnor2_1 _11654_ (.Y(_05660_),
    .A(net874),
    .B(net584));
 sg13g2_nor2_1 _11655_ (.A(net587),
    .B(_05660_),
    .Y(_05661_));
 sg13g2_a221oi_1 _11656_ (.B2(net647),
    .C1(_05661_),
    .B1(_05659_),
    .A1(net594),
    .Y(_05662_),
    .A2(_05653_));
 sg13g2_buf_2 fanout611 (.A(_05276_),
    .X(net611));
 sg13g2_o21ai_1 _11658_ (.B1(_05436_),
    .Y(_05664_),
    .A1(net912),
    .A2(_05573_));
 sg13g2_a22oi_1 _11659_ (.Y(_05665_),
    .B1(_05662_),
    .B2(_05664_),
    .A2(_05598_),
    .A1(_05585_));
 sg13g2_buf_1 fanout610 (.A(_05288_),
    .X(net610));
 sg13g2_or3_1 _11661_ (.A(_05433_),
    .B(_05566_),
    .C(_05665_),
    .X(_05667_));
 sg13g2_nand4_1 _11662_ (.B(_05243_),
    .C(_05432_),
    .A(_04790_),
    .Y(_05668_),
    .D(_05667_));
 sg13g2_nand2_1 _11663_ (.Y(_05669_),
    .A(_05232_),
    .B(_05668_));
 sg13g2_buf_1 fanout609 (.A(net610),
    .X(net609));
 sg13g2_xor2_1 _11665_ (.B(_04110_),
    .A(net633),
    .X(_05671_));
 sg13g2_buf_2 fanout608 (.A(net610),
    .X(net608));
 sg13g2_nor2_2 _11667_ (.A(_04025_),
    .B(_04049_),
    .Y(_05673_));
 sg13g2_buf_2 fanout607 (.A(net610),
    .X(net607));
 sg13g2_xnor2_1 _11669_ (.Y(_05675_),
    .A(_05673_),
    .B(_04060_));
 sg13g2_nand2b_1 _11670_ (.Y(_05676_),
    .B(_05675_),
    .A_N(_05671_));
 sg13g2_xnor2_1 _11671_ (.Y(_05677_),
    .A(net631),
    .B(_04173_));
 sg13g2_xnor2_1 _11672_ (.Y(_05678_),
    .A(_03901_),
    .B(_04177_));
 sg13g2_buf_2 fanout606 (.A(net607),
    .X(net606));
 sg13g2_nor3_2 _11674_ (.A(_05676_),
    .B(_05677_),
    .C(_05678_),
    .Y(_05680_));
 sg13g2_buf_2 fanout605 (.A(net607),
    .X(net605));
 sg13g2_and3_1 _11676_ (.X(_05682_),
    .A(net338),
    .B(_05680_),
    .C(_04400_));
 sg13g2_buf_1 fanout604 (.A(_05316_),
    .X(net604));
 sg13g2_a21o_2 _11678_ (.A2(_04372_),
    .A1(_04368_),
    .B1(_04388_),
    .X(_05684_));
 sg13g2_buf_2 fanout603 (.A(_05316_),
    .X(net603));
 sg13g2_and2_1 _11680_ (.A(_04278_),
    .B(_04285_),
    .X(_05686_));
 sg13g2_buf_2 fanout602 (.A(_05411_),
    .X(net602));
 sg13g2_and2_1 _11682_ (.A(_04191_),
    .B(_05686_),
    .X(_05688_));
 sg13g2_a21oi_1 _11683_ (.A1(_04278_),
    .A2(_04285_),
    .Y(_05689_),
    .B1(_04191_));
 sg13g2_nor2_1 _11684_ (.A(_05689_),
    .B(_04235_),
    .Y(_05690_));
 sg13g2_a22oi_1 _11685_ (.Y(_05691_),
    .B1(_05688_),
    .B2(_05690_),
    .A2(_04396_),
    .A1(_05684_));
 sg13g2_nand2b_1 _11686_ (.Y(_05692_),
    .B(_04389_),
    .A_N(_04396_));
 sg13g2_buf_1 fanout601 (.A(_05420_),
    .X(net601));
 sg13g2_nor2b_1 _11688_ (.A(_05691_),
    .B_N(_05692_),
    .Y(_05694_));
 sg13g2_xnor2_1 _11689_ (.Y(_05695_),
    .A(net872),
    .B(_04347_));
 sg13g2_nand2_1 _11690_ (.Y(_05696_),
    .A(_05694_),
    .B(_05695_));
 sg13g2_nor2_1 _11691_ (.A(_05694_),
    .B(_05695_),
    .Y(_05697_));
 sg13g2_inv_1 _11692_ (.Y(_05698_),
    .A(_04350_));
 sg13g2_a22oi_1 _11693_ (.Y(_05699_),
    .B1(_05697_),
    .B2(_05698_),
    .A2(_05696_),
    .A1(net630));
 sg13g2_nor2_1 _11694_ (.A(net629),
    .B(_04352_),
    .Y(_05700_));
 sg13g2_a22oi_1 _11695_ (.Y(_05701_),
    .B1(_05700_),
    .B2(_04350_),
    .A2(_04353_),
    .A1(_05692_));
 sg13g2_or3_1 _11696_ (.A(net635),
    .B(_05699_),
    .C(_05701_),
    .X(_05702_));
 sg13g2_a22oi_1 _11697_ (.Y(_05703_),
    .B1(_05682_),
    .B2(_05702_),
    .A2(_04400_),
    .A1(_04183_));
 sg13g2_nand2b_1 _11698_ (.Y(_05704_),
    .B(_05680_),
    .A_N(_04289_));
 sg13g2_a21oi_1 _11699_ (.A1(_05232_),
    .A2(_05668_),
    .Y(_05705_),
    .B1(_05704_));
 sg13g2_nor4_1 _11700_ (.A(_05694_),
    .B(_03887_),
    .C(_04350_),
    .D(_05700_),
    .Y(_05706_));
 sg13g2_nand2b_1 _11701_ (.Y(_05707_),
    .B(_04183_),
    .A_N(_04289_));
 sg13g2_nand2_1 _11702_ (.Y(_05708_),
    .A(_05706_),
    .B(_05707_));
 sg13g2_nor3_1 _11703_ (.A(net1240),
    .B(_03881_),
    .C(_03865_),
    .Y(_05709_));
 sg13g2_buf_2 fanout600 (.A(net601),
    .X(net600));
 sg13g2_buf_2 fanout599 (.A(_05427_),
    .X(net599));
 sg13g2_buf_2 fanout598 (.A(_05495_),
    .X(net598));
 sg13g2_buf_2 fanout597 (.A(net598),
    .X(net597));
 sg13g2_buf_2 fanout596 (.A(_05563_),
    .X(net596));
 sg13g2_buf_2 fanout595 (.A(_05599_),
    .X(net595));
 sg13g2_buf_2 fanout594 (.A(net595),
    .X(net594));
 sg13g2_buf_2 fanout593 (.A(net595),
    .X(net593));
 sg13g2_buf_2 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_2 fanout591 (.A(net592),
    .X(net591));
 sg13g2_mux4_1 _11714_ (.S0(net639),
    .A0(net621),
    .A1(_04685_),
    .A2(_05225_),
    .A3(_05223_),
    .S1(net578),
    .X(_05720_));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(_05599_));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(net590));
 sg13g2_buf_2 fanout588 (.A(net589),
    .X(net588));
 sg13g2_mux2_1 _11718_ (.A0(net625),
    .A1(_04550_),
    .S(net581),
    .X(_05724_));
 sg13g2_buf_2 fanout587 (.A(_05639_),
    .X(net587));
 sg13g2_mux2_1 _11720_ (.A0(_05198_),
    .A1(net623),
    .S(net571),
    .X(_05726_));
 sg13g2_mux2_1 _11721_ (.A0(_05724_),
    .A1(_05726_),
    .S(net642),
    .X(_05727_));
 sg13g2_nor2_1 _11722_ (.A(net383),
    .B(_05727_),
    .Y(_05728_));
 sg13g2_a21oi_1 _11723_ (.A1(net383),
    .A2(_05720_),
    .Y(_05729_),
    .B1(_05728_));
 sg13g2_buf_1 fanout586 (.A(_05650_),
    .X(net586));
 sg13g2_buf_1 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_2 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_2 fanout583 (.A(net585),
    .X(net583));
 sg13g2_mux4_1 _11728_ (.S0(net588),
    .A0(_03989_),
    .A1(net631),
    .A2(net632),
    .A3(net568),
    .S1(net579),
    .X(_05734_));
 sg13g2_nor2_2 _11729_ (.A(_04261_),
    .B(_04276_),
    .Y(_05735_));
 sg13g2_mux2_1 _11730_ (.A0(net626),
    .A1(_05735_),
    .S(net579),
    .X(_05736_));
 sg13g2_mux2_1 _11731_ (.A0(_04235_),
    .A1(net628),
    .S(net570),
    .X(_05737_));
 sg13g2_mux2_1 _11732_ (.A0(_05736_),
    .A1(_05737_),
    .S(net641),
    .X(_05738_));
 sg13g2_mux2_1 _11733_ (.A0(_05734_),
    .A1(_05738_),
    .S(net383),
    .X(_05739_));
 sg13g2_or2_1 _11734_ (.X(_05740_),
    .B(_05739_),
    .A(net364));
 sg13g2_o21ai_1 _11735_ (.B1(_05740_),
    .Y(_05741_),
    .A1(net395),
    .A2(_05729_));
 sg13g2_buf_2 fanout582 (.A(net585),
    .X(net582));
 sg13g2_buf_2 fanout581 (.A(net586),
    .X(net581));
 sg13g2_buf_2 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579));
 sg13g2_and2_1 _11740_ (.A(net617),
    .B(net582),
    .X(_05746_));
 sg13g2_buf_2 fanout578 (.A(net581),
    .X(net578));
 sg13g2_a21o_1 _11742_ (.A2(net573),
    .A1(net618),
    .B1(_05746_),
    .X(_05748_));
 sg13g2_mux2_1 _11743_ (.A0(_05177_),
    .A1(_04928_),
    .S(net586),
    .X(_05749_));
 sg13g2_mux2_1 _11744_ (.A0(_05748_),
    .A1(_05749_),
    .S(net646),
    .X(_05750_));
 sg13g2_buf_1 fanout577 (.A(_05654_),
    .X(net577));
 sg13g2_buf_1 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_1 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_2 fanout574 (.A(net575),
    .X(net574));
 sg13g2_nor2_1 _11749_ (.A(net613),
    .B(net574),
    .Y(_05755_));
 sg13g2_a21oi_1 _11750_ (.A1(net402),
    .A2(net574),
    .Y(_05756_),
    .B1(_05755_));
 sg13g2_nand3_1 _11751_ (.B(_05104_),
    .C(_05118_),
    .A(_05095_),
    .Y(_05757_));
 sg13g2_buf_2 fanout573 (.A(net575),
    .X(net573));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(net573));
 sg13g2_nor2_1 _11754_ (.A(net566),
    .B(net575),
    .Y(_05760_));
 sg13g2_a22oi_1 _11755_ (.Y(_05761_),
    .B1(_05760_),
    .B2(net595),
    .A2(net574),
    .A1(net401));
 sg13g2_a22oi_1 _11756_ (.Y(_05762_),
    .B1(_05761_),
    .B2(net388),
    .A2(_05756_),
    .A1(net594));
 sg13g2_a21oi_1 _11757_ (.A1(net388),
    .A2(_05750_),
    .Y(_05763_),
    .B1(_05762_));
 sg13g2_buf_2 fanout571 (.A(net577),
    .X(net571));
 sg13g2_buf_2 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_2 fanout569 (.A(net571),
    .X(net569));
 sg13g2_nor2_1 _11761_ (.A(net591),
    .B(net600),
    .Y(_05767_));
 sg13g2_a21oi_1 _11762_ (.A1(net591),
    .A2(net599),
    .Y(_05768_),
    .B1(_05767_));
 sg13g2_buf_2 fanout568 (.A(_05673_),
    .X(net568));
 sg13g2_nor2_1 _11764_ (.A(net591),
    .B(net603),
    .Y(_05770_));
 sg13g2_a22oi_1 _11765_ (.Y(_05771_),
    .B1(net572),
    .B2(_05770_),
    .A2(net611),
    .A1(net591));
 sg13g2_a21oi_1 _11766_ (.A1(net572),
    .A2(_05768_),
    .Y(_05772_),
    .B1(_05771_));
 sg13g2_nor2_1 _11767_ (.A(net587),
    .B(net574),
    .Y(_05773_));
 sg13g2_a22oi_1 _11768_ (.Y(_05774_),
    .B1(_05773_),
    .B2(net594),
    .A2(net574),
    .A1(net391));
 sg13g2_buf_1 fanout567 (.A(_05757_),
    .X(net567));
 sg13g2_nand4_1 _11770_ (.B(_05578_),
    .C(_05580_),
    .A(net912),
    .Y(_05776_),
    .D(_05582_));
 sg13g2_buf_2 fanout566 (.A(_05757_),
    .X(net566));
 sg13g2_nor2_1 _11772_ (.A(_05776_),
    .B(net585),
    .Y(_05778_));
 sg13g2_a22oi_1 _11773_ (.Y(_05779_),
    .B1(_05778_),
    .B2(net644),
    .A2(net585),
    .A1(net647));
 sg13g2_nor3_1 _11774_ (.A(net389),
    .B(_05774_),
    .C(_05779_),
    .Y(_05780_));
 sg13g2_a22oi_1 _11775_ (.Y(_05781_),
    .B1(_05780_),
    .B2(net400),
    .A2(_05772_),
    .A1(net389));
 sg13g2_a22oi_1 _11776_ (.Y(_05782_),
    .B1(_05781_),
    .B2(net608),
    .A2(_05763_),
    .A1(net399));
 sg13g2_a21o_1 _11777_ (.A2(_05741_),
    .A1(net606),
    .B1(_05782_),
    .X(_05783_));
 sg13g2_nor2_1 _11778_ (.A(net983),
    .B(_03865_),
    .Y(_05784_));
 sg13g2_nand3_1 _11779_ (.B(_03861_),
    .C(_05784_),
    .A(net934),
    .Y(_05785_));
 sg13g2_buf_1 fanout565 (.A(_05798_),
    .X(net565));
 sg13g2_buf_2 fanout564 (.A(net565),
    .X(net564));
 sg13g2_nor2_1 _11782_ (.A(net608),
    .B(net869),
    .Y(_05788_));
 sg13g2_buf_2 fanout563 (.A(_07398_),
    .X(net563));
 sg13g2_inv_1 _11784_ (.Y(_05790_),
    .A(net358));
 sg13g2_nand3_1 _11785_ (.B(net590),
    .C(net581),
    .A(net648),
    .Y(_05791_));
 sg13g2_buf_2 fanout562 (.A(_07398_),
    .X(net562));
 sg13g2_nand2_1 _11787_ (.Y(_05793_),
    .A(net369),
    .B(net359));
 sg13g2_buf_1 fanout561 (.A(_07492_),
    .X(net561));
 sg13g2_nor4_1 _11789_ (.A(net835),
    .B(_05790_),
    .C(_05791_),
    .D(_05793_),
    .Y(_05795_));
 sg13g2_buf_2 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_2 fanout559 (.A(net561),
    .X(net559));
 sg13g2_nand3_1 _11792_ (.B(_03864_),
    .C(_03876_),
    .A(_03857_),
    .Y(_05798_));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_nand2_1 _11794_ (.Y(_05800_),
    .A(net845),
    .B(net564));
 sg13g2_buf_2 fanout557 (.A(_07569_),
    .X(net557));
 sg13g2_buf_2 fanout556 (.A(net557),
    .X(net556));
 sg13g2_xnor2_1 _11797_ (.Y(_05803_),
    .A(net648),
    .B(net642));
 sg13g2_and3_1 _11798_ (.X(_05804_),
    .A(net934),
    .B(_03861_),
    .C(_05784_));
 sg13g2_buf_2 fanout555 (.A(_07748_),
    .X(net555));
 sg13g2_a22oi_1 _11800_ (.Y(_05806_),
    .B1(_05803_),
    .B2(net831),
    .A2(net356),
    .A1(net848));
 sg13g2_a22oi_1 _11801_ (.Y(_05807_),
    .B1(_05795_),
    .B2(_05806_),
    .A2(_05783_),
    .A1(net869));
 sg13g2_o21ai_1 _11802_ (.B1(_05807_),
    .Y(_05808_),
    .A1(_05705_),
    .A2(_05708_));
 sg13g2_inv_1 _11803_ (.Y(_05809_),
    .A(_05808_));
 sg13g2_o21ai_1 _11804_ (.B1(_05809_),
    .Y(net66),
    .A1(_03887_),
    .A2(_05703_));
 sg13g2_nand2b_1 _11805_ (.Y(_05810_),
    .B(_03865_),
    .A_N(net1249));
 sg13g2_buf_2 fanout554 (.A(net555),
    .X(net554));
 sg13g2_inv_1 _11807_ (.Y(net98),
    .A(net863));
 sg13g2_buf_2 fanout553 (.A(net555),
    .X(net553));
 sg13g2_buf_2 fanout552 (.A(net555),
    .X(net552));
 sg13g2_nand2_1 _11810_ (.Y(_05814_),
    .A(net1237),
    .B(_05784_));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout550 (.A(_07748_),
    .X(net550));
 sg13g2_buf_2 fanout549 (.A(net550),
    .X(net549));
 sg13g2_nor2_1 _11814_ (.A(net385),
    .B(net397),
    .Y(_05818_));
 sg13g2_buf_2 fanout548 (.A(net550),
    .X(net548));
 sg13g2_nand2_1 _11816_ (.Y(_05820_),
    .A(net647),
    .B(net645));
 sg13g2_nand2b_1 _11817_ (.Y(_05821_),
    .B(net594),
    .A_N(net587));
 sg13g2_a21oi_1 _11818_ (.A1(_05820_),
    .A2(_05821_),
    .Y(_05822_),
    .B1(net574));
 sg13g2_and2_1 _11819_ (.A(_05818_),
    .B(_05822_),
    .X(_05823_));
 sg13g2_buf_1 fanout547 (.A(net550),
    .X(net547));
 sg13g2_buf_2 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_1 fanout545 (.A(_07792_),
    .X(net545));
 sg13g2_buf_2 fanout544 (.A(_07792_),
    .X(net544));
 sg13g2_a21o_1 _11824_ (.A2(net574),
    .A1(net401),
    .B1(_05760_),
    .X(_05828_));
 sg13g2_nand3_1 _11825_ (.B(_05058_),
    .C(_05083_),
    .A(net912),
    .Y(_05829_));
 sg13g2_buf_1 fanout543 (.A(_07797_),
    .X(net543));
 sg13g2_buf_1 fanout542 (.A(net543),
    .X(net542));
 sg13g2_nor2_1 _11828_ (.A(net617),
    .B(net582),
    .Y(_05832_));
 sg13g2_a21oi_1 _11829_ (.A1(net354),
    .A2(net582),
    .Y(_05833_),
    .B1(_05832_));
 sg13g2_mux2_1 _11830_ (.A0(_05828_),
    .A1(_05833_),
    .S(net643),
    .X(_05834_));
 sg13g2_and3_2 _11831_ (.X(_05835_),
    .A(_04517_),
    .B(_04528_),
    .C(_04548_));
 sg13g2_buf_2 fanout541 (.A(net542),
    .X(net541));
 sg13g2_mux2_1 _11833_ (.A0(_05835_),
    .A1(net618),
    .S(net586),
    .X(_05837_));
 sg13g2_mux2_1 _11834_ (.A0(_05749_),
    .A1(_05837_),
    .S(net646),
    .X(_05838_));
 sg13g2_and2_1 _11835_ (.A(net387),
    .B(_05838_),
    .X(_05839_));
 sg13g2_a21oi_1 _11836_ (.A1(net376),
    .A2(_05834_),
    .Y(_05840_),
    .B1(_05839_));
 sg13g2_buf_2 fanout540 (.A(net543),
    .X(net540));
 sg13g2_and2_1 _11838_ (.A(net912),
    .B(_05656_),
    .X(_05842_));
 sg13g2_buf_2 fanout539 (.A(net543),
    .X(net539));
 sg13g2_mux4_1 _11840_ (.S0(net583),
    .A0(net611),
    .A1(net596),
    .A2(net391),
    .A3(_05842_),
    .S1(net592),
    .X(_05844_));
 sg13g2_buf_2 fanout538 (.A(net543),
    .X(net538));
 sg13g2_buf_2 fanout537 (.A(net538),
    .X(net537));
 sg13g2_mux4_1 _11843_ (.S0(net583),
    .A0(net613),
    .A1(net602),
    .A2(net600),
    .A3(net603),
    .S1(net592),
    .X(_05847_));
 sg13g2_nor2_1 _11844_ (.A(net376),
    .B(_05847_),
    .Y(_05848_));
 sg13g2_a22oi_1 _11845_ (.Y(_05849_),
    .B1(_05848_),
    .B2(net400),
    .A2(_05844_),
    .A1(net375));
 sg13g2_a22oi_1 _11846_ (.Y(_05850_),
    .B1(_05849_),
    .B2(net824),
    .A2(_05840_),
    .A1(net400));
 sg13g2_buf_1 fanout536 (.A(net537),
    .X(net536));
 sg13g2_a22oi_1 _11848_ (.Y(_05852_),
    .B1(_05850_),
    .B2(net608),
    .A2(_05823_),
    .A1(net824));
 sg13g2_nor2_1 _11849_ (.A(_04391_),
    .B(net825),
    .Y(_05853_));
 sg13g2_buf_2 fanout535 (.A(net537),
    .X(net535));
 sg13g2_nand2_1 _11851_ (.Y(_05855_),
    .A(net620),
    .B(net571));
 sg13g2_o21ai_1 _11852_ (.B1(_05855_),
    .Y(_05856_),
    .A1(_04502_),
    .A2(net571));
 sg13g2_mux2_1 _11853_ (.A0(_05726_),
    .A1(_05856_),
    .S(net642),
    .X(_05857_));
 sg13g2_mux2_1 _11854_ (.A0(net621),
    .A1(_05223_),
    .S(net590),
    .X(_05858_));
 sg13g2_mux2_1 _11855_ (.A0(_04050_),
    .A1(_04685_),
    .S(net590),
    .X(_05859_));
 sg13g2_mux2_1 _11856_ (.A0(_05858_),
    .A1(_05859_),
    .S(net570),
    .X(_05860_));
 sg13g2_nor2_1 _11857_ (.A(net370),
    .B(_05860_),
    .Y(_05861_));
 sg13g2_a21oi_1 _11858_ (.A1(net374),
    .A2(_05857_),
    .Y(_05862_),
    .B1(_05861_));
 sg13g2_nand2_1 _11859_ (.Y(_05863_),
    .A(net364),
    .B(_05862_));
 sg13g2_mux4_1 _11860_ (.S0(net590),
    .A0(_05735_),
    .A1(_03989_),
    .A2(_04166_),
    .A3(net632),
    .S1(net580),
    .X(_05864_));
 sg13g2_and2_1 _11861_ (.A(net370),
    .B(_05864_),
    .X(_05865_));
 sg13g2_nand2b_1 _11862_ (.Y(_05866_),
    .B(net570),
    .A_N(net627));
 sg13g2_inv_1 _11863_ (.Y(_05867_),
    .A(_05866_));
 sg13g2_or2_2 _11864_ (.X(_05868_),
    .B(_04233_),
    .A(_04211_));
 sg13g2_buf_1 fanout534 (.A(_07882_),
    .X(net534));
 sg13g2_nor2_1 _11866_ (.A(_05868_),
    .B(net641),
    .Y(_05870_));
 sg13g2_a22oi_1 _11867_ (.Y(_05871_),
    .B1(net570),
    .B2(_05870_),
    .A2(net641),
    .A1(net626));
 sg13g2_buf_2 fanout533 (.A(net534),
    .X(net533));
 sg13g2_nor3_1 _11869_ (.A(net370),
    .B(_05867_),
    .C(_05871_),
    .Y(_05873_));
 sg13g2_or3_1 _11870_ (.A(net361),
    .B(_05865_),
    .C(_05873_),
    .X(_05874_));
 sg13g2_nand2_1 _11871_ (.Y(_05875_),
    .A(_05863_),
    .B(_05874_));
 sg13g2_a21o_2 _11872_ (.A2(_05282_),
    .A1(_05280_),
    .B1(_05287_),
    .X(_05876_));
 sg13g2_buf_2 fanout532 (.A(net533),
    .X(net532));
 sg13g2_nor2_1 _11874_ (.A(net911),
    .B(_05876_),
    .Y(_05878_));
 sg13g2_a21oi_1 _11875_ (.A1(net159),
    .A2(net911),
    .Y(_05879_),
    .B1(_05878_));
 sg13g2_buf_2 fanout531 (.A(net533),
    .X(net531));
 sg13g2_buf_2 fanout530 (.A(net533),
    .X(net530));
 sg13g2_buf_2 fanout529 (.A(net533),
    .X(net529));
 sg13g2_a21oi_1 _11879_ (.A1(_05684_),
    .A2(net580),
    .Y(_05883_),
    .B1(net589));
 sg13g2_a21o_1 _11880_ (.A2(_05737_),
    .A1(net589),
    .B1(_05883_),
    .X(_05884_));
 sg13g2_buf_2 fanout528 (.A(net534),
    .X(net528));
 sg13g2_a21oi_1 _11882_ (.A1(net381),
    .A2(_05884_),
    .Y(_05886_),
    .B1(_05865_));
 sg13g2_nand2_1 _11883_ (.Y(_05887_),
    .A(net397),
    .B(_05886_));
 sg13g2_nand2_2 _11884_ (.Y(_05888_),
    .A(_04391_),
    .B(net868));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_a21oi_1 _11886_ (.A1(_05863_),
    .A2(_05887_),
    .Y(_05890_),
    .B1(_05888_));
 sg13g2_a22oi_1 _11887_ (.Y(_05891_),
    .B1(net350),
    .B2(_05890_),
    .A2(_05875_),
    .A1(_05853_));
 sg13g2_buf_2 fanout526 (.A(net528),
    .X(net526));
 sg13g2_buf_2 fanout525 (.A(_07926_),
    .X(net525));
 sg13g2_o21ai_1 _11890_ (.B1(net834),
    .Y(_05894_),
    .A1(_05852_),
    .A2(_05891_));
 sg13g2_buf_2 fanout524 (.A(net525),
    .X(net524));
 sg13g2_xnor2_1 _11892_ (.Y(_05896_),
    .A(net587),
    .B(_05660_));
 sg13g2_o21ai_1 _11893_ (.B1(_05820_),
    .Y(_05897_),
    .A1(net876),
    .A2(net645));
 sg13g2_xor2_1 _11894_ (.B(_05897_),
    .A(_05896_),
    .X(_05898_));
 sg13g2_buf_1 fanout523 (.A(_07968_),
    .X(net523));
 sg13g2_buf_2 fanout522 (.A(net523),
    .X(net522));
 sg13g2_buf_2 fanout521 (.A(net523),
    .X(net521));
 sg13g2_and3_1 _11898_ (.X(_05902_),
    .A(net1238),
    .B(_02576_),
    .C(_03851_));
 sg13g2_buf_2 fanout520 (.A(net521),
    .X(net520));
 sg13g2_buf_2 fanout519 (.A(net521),
    .X(net519));
 sg13g2_o21ai_1 _11901_ (.B1(net845),
    .Y(_05905_),
    .A1(net820),
    .A2(net587));
 sg13g2_nand2b_1 _11902_ (.Y(_05906_),
    .B(_05905_),
    .A_N(_05660_));
 sg13g2_o21ai_1 _11903_ (.B1(_05906_),
    .Y(_05907_),
    .A1(net845),
    .A2(net587));
 sg13g2_buf_2 fanout518 (.A(net521),
    .X(net518));
 sg13g2_nor2_1 _11905_ (.A(net850),
    .B(_05896_),
    .Y(_05909_));
 sg13g2_a22oi_1 _11906_ (.Y(_05910_),
    .B1(_05909_),
    .B2(net833),
    .A2(_05907_),
    .A1(net636));
 sg13g2_o21ai_1 _11907_ (.B1(_05910_),
    .Y(_05911_),
    .A1(net357),
    .A2(_05898_));
 sg13g2_and2_1 _11908_ (.A(_05894_),
    .B(_05911_),
    .X(net77));
 sg13g2_nand2_2 _11909_ (.Y(_05912_),
    .A(net351),
    .B(net869));
 sg13g2_buf_2 fanout517 (.A(_07968_),
    .X(net517));
 sg13g2_inv_1 _11911_ (.Y(_05914_),
    .A(_05912_));
 sg13g2_buf_2 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_2 fanout515 (.A(net517),
    .X(net515));
 sg13g2_nand2_2 _11914_ (.Y(_05917_),
    .A(_05128_),
    .B(_05162_));
 sg13g2_nor2_1 _11915_ (.A(_04928_),
    .B(net582),
    .Y(_05918_));
 sg13g2_a21oi_1 _11916_ (.A1(_05917_),
    .A2(net582),
    .Y(_05919_),
    .B1(_05918_));
 sg13g2_mux2_1 _11917_ (.A0(_05833_),
    .A1(_05919_),
    .S(net643),
    .X(_05920_));
 sg13g2_nand2_1 _11918_ (.Y(_05921_),
    .A(_04830_),
    .B(net581));
 sg13g2_nand2_1 _11919_ (.Y(_05922_),
    .A(_05198_),
    .B(net571));
 sg13g2_and2_1 _11920_ (.A(_05921_),
    .B(_05922_),
    .X(_05923_));
 sg13g2_mux2_1 _11921_ (.A0(_05837_),
    .A1(_05923_),
    .S(net646),
    .X(_05924_));
 sg13g2_mux2_1 _11922_ (.A0(_05920_),
    .A1(_05924_),
    .S(net387),
    .X(_05925_));
 sg13g2_nand2_1 _11923_ (.Y(_05926_),
    .A(net912),
    .B(net597));
 sg13g2_mux4_1 _11924_ (.S0(net644),
    .A0(_05434_),
    .A1(net603),
    .A2(_05776_),
    .A3(_05926_),
    .S1(net584),
    .X(_05927_));
 sg13g2_nor2_1 _11925_ (.A(net591),
    .B(net566),
    .Y(_05928_));
 sg13g2_a21oi_1 _11926_ (.A1(net591),
    .A2(_05237_),
    .Y(_05929_),
    .B1(_05928_));
 sg13g2_mux2_1 _11927_ (.A0(_05768_),
    .A1(_05929_),
    .S(net572),
    .X(_05930_));
 sg13g2_mux2_1 _11928_ (.A0(_05927_),
    .A1(_05930_),
    .S(net389),
    .X(_05931_));
 sg13g2_nand2_1 _11929_ (.Y(_05932_),
    .A(net368),
    .B(_05931_));
 sg13g2_o21ai_1 _11930_ (.B1(_05932_),
    .Y(_05933_),
    .A1(net366),
    .A2(_05925_));
 sg13g2_mux2_1 _11931_ (.A0(net647),
    .A1(net596),
    .S(net583),
    .X(_05934_));
 sg13g2_nor3_1 _11932_ (.A(net592),
    .B(net587),
    .C(net572),
    .Y(_05935_));
 sg13g2_a21o_1 _11933_ (.A2(_05934_),
    .A1(net592),
    .B1(_05935_),
    .X(_05936_));
 sg13g2_buf_2 fanout514 (.A(net515),
    .X(net514));
 sg13g2_nand2_1 _11935_ (.Y(_05938_),
    .A(_05818_),
    .B(_05936_));
 sg13g2_mux2_1 _11936_ (.A0(net626),
    .A1(net627),
    .S(net640),
    .X(_05939_));
 sg13g2_nand2b_1 _11937_ (.Y(_05940_),
    .B(net579),
    .A_N(_05939_));
 sg13g2_buf_1 fanout513 (.A(_08067_),
    .X(net513));
 sg13g2_a21o_2 _11939_ (.A2(_04142_),
    .A1(_04121_),
    .B1(_04165_),
    .X(_05942_));
 sg13g2_buf_2 fanout512 (.A(_08067_),
    .X(net512));
 sg13g2_mux4_1 _11941_ (.S0(net639),
    .A0(_04278_),
    .A1(_05868_),
    .A2(_05942_),
    .A3(_04177_),
    .S1(net579),
    .X(_05944_));
 sg13g2_buf_2 fanout511 (.A(_08091_),
    .X(net511));
 sg13g2_nand2_1 _11943_ (.Y(_05946_),
    .A(net370),
    .B(_05944_));
 sg13g2_o21ai_1 _11944_ (.B1(_05946_),
    .Y(_05947_),
    .A1(net370),
    .A2(_05940_));
 sg13g2_mux4_1 _11945_ (.S0(net642),
    .A0(net624),
    .A1(net623),
    .A2(net620),
    .A3(_04725_),
    .S1(net577),
    .X(_05948_));
 sg13g2_and2_1 _11946_ (.A(_04617_),
    .B(_04631_),
    .X(_05949_));
 sg13g2_buf_2 fanout510 (.A(net511),
    .X(net510));
 sg13g2_mux4_1 _11948_ (.S0(net589),
    .A0(net632),
    .A1(net568),
    .A2(_05215_),
    .A3(_05949_),
    .S1(net579),
    .X(_05951_));
 sg13g2_mux2_1 _11949_ (.A0(_05948_),
    .A1(_05951_),
    .S(net384),
    .X(_05952_));
 sg13g2_nor2_1 _11950_ (.A(net397),
    .B(_05952_),
    .Y(_05953_));
 sg13g2_a21oi_1 _11951_ (.A1(net398),
    .A2(_05947_),
    .Y(_05954_),
    .B1(_05953_));
 sg13g2_nor2_1 _11952_ (.A(_05888_),
    .B(_05954_),
    .Y(_05955_));
 sg13g2_nand2_2 _11953_ (.Y(_05956_),
    .A(net1253),
    .B(net870));
 sg13g2_buf_1 fanout509 (.A(_08130_),
    .X(net509));
 sg13g2_nand2_1 _11955_ (.Y(_05958_),
    .A(_05866_),
    .B(_05940_));
 sg13g2_nor2_1 _11956_ (.A(net392),
    .B(_05951_),
    .Y(_05959_));
 sg13g2_a22oi_1 _11957_ (.Y(_05960_),
    .B1(_05959_),
    .B2(net370),
    .A2(_05958_),
    .A1(net394));
 sg13g2_nor2_1 _11958_ (.A(net393),
    .B(_05948_),
    .Y(_05961_));
 sg13g2_a22oi_1 _11959_ (.Y(_05962_),
    .B1(_05961_),
    .B2(net382),
    .A2(_05944_),
    .A1(net394));
 sg13g2_nor3_1 _11960_ (.A(_05956_),
    .B(_05960_),
    .C(_05962_),
    .Y(_05963_));
 sg13g2_nor3_1 _11961_ (.A(net352),
    .B(_05955_),
    .C(_05963_),
    .Y(_05964_));
 sg13g2_a221oi_1 _11962_ (.B2(_05788_),
    .C1(_05964_),
    .B1(_05938_),
    .A1(_05914_),
    .Y(_05965_),
    .A2(_05933_));
 sg13g2_buf_2 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_1 fanout507 (.A(net509),
    .X(net507));
 sg13g2_buf_2 fanout506 (.A(net507),
    .X(net506));
 sg13g2_xnor2_1 _11966_ (.Y(_05969_),
    .A(net874),
    .B(net389));
 sg13g2_xnor2_1 _11967_ (.Y(_05970_),
    .A(_05776_),
    .B(_05969_));
 sg13g2_nor2_1 _11968_ (.A(net596),
    .B(_05969_),
    .Y(_05971_));
 sg13g2_nand3_1 _11969_ (.B(net596),
    .C(_05969_),
    .A(net850),
    .Y(_05972_));
 sg13g2_o21ai_1 _11970_ (.B1(_05972_),
    .Y(_05973_),
    .A1(net845),
    .A2(_05971_));
 sg13g2_xor2_1 _11971_ (.B(_05970_),
    .A(_05662_),
    .X(_05974_));
 sg13g2_nor2_1 _11972_ (.A(net357),
    .B(_05974_),
    .Y(_05975_));
 sg13g2_a221oi_1 _11973_ (.B2(net636),
    .C1(_05975_),
    .B1(_05973_),
    .A1(net820),
    .Y(_05976_),
    .A2(_05970_));
 sg13g2_nor2_1 _11974_ (.A(net833),
    .B(_05976_),
    .Y(_05977_));
 sg13g2_a21o_1 _11975_ (.A2(_05965_),
    .A1(net833),
    .B1(_05977_),
    .X(net88));
 sg13g2_buf_2 fanout505 (.A(net507),
    .X(net505));
 sg13g2_nor2_1 _11977_ (.A(net590),
    .B(_05724_),
    .Y(_05979_));
 sg13g2_a21oi_1 _11978_ (.A1(net590),
    .A2(_05923_),
    .Y(_05980_),
    .B1(_05979_));
 sg13g2_mux2_1 _11979_ (.A0(_05748_),
    .A1(_05919_),
    .S(net593),
    .X(_05981_));
 sg13g2_nor2_1 _11980_ (.A(net388),
    .B(_05981_),
    .Y(_05982_));
 sg13g2_a21oi_1 _11981_ (.A1(net388),
    .A2(_05980_),
    .Y(_05983_),
    .B1(_05982_));
 sg13g2_nor2_1 _11982_ (.A(net566),
    .B(net584),
    .Y(_05984_));
 sg13g2_a21oi_1 _11983_ (.A1(_05362_),
    .A2(net584),
    .Y(_05985_),
    .B1(_05984_));
 sg13g2_mux2_1 _11984_ (.A0(_05756_),
    .A1(_05985_),
    .S(net594),
    .X(_05986_));
 sg13g2_nor2_1 _11985_ (.A(net644),
    .B(net604),
    .Y(_05987_));
 sg13g2_a22oi_1 _11986_ (.Y(_05988_),
    .B1(net584),
    .B2(_05987_),
    .A2(net599),
    .A1(net643));
 sg13g2_nor2_1 _11987_ (.A(net643),
    .B(_05926_),
    .Y(_05989_));
 sg13g2_a22oi_1 _11988_ (.Y(_05990_),
    .B1(net574),
    .B2(_05989_),
    .A2(net611),
    .A1(net643));
 sg13g2_or3_1 _11989_ (.A(net390),
    .B(_05988_),
    .C(_05990_),
    .X(_05991_));
 sg13g2_o21ai_1 _11990_ (.B1(_05991_),
    .Y(_05992_),
    .A1(net376),
    .A2(_05986_));
 sg13g2_mux2_1 _11991_ (.A0(_05983_),
    .A1(_05992_),
    .S(net366),
    .X(_05993_));
 sg13g2_mux4_1 _11992_ (.S0(net570),
    .A0(net612),
    .A1(_05223_),
    .A2(_05225_),
    .A3(net621),
    .S1(net641),
    .X(_05994_));
 sg13g2_mux4_1 _11993_ (.S0(net589),
    .A0(net631),
    .A1(net632),
    .A2(net568),
    .A3(_05215_),
    .S1(net580),
    .X(_05995_));
 sg13g2_nor2_1 _11994_ (.A(net378),
    .B(_05995_),
    .Y(_05996_));
 sg13g2_a21oi_1 _11995_ (.A1(net374),
    .A2(_05994_),
    .Y(_05997_),
    .B1(_05996_));
 sg13g2_nor2_1 _11996_ (.A(net397),
    .B(_05997_),
    .Y(_05998_));
 sg13g2_or3_1 _11997_ (.A(net642),
    .B(net628),
    .C(net577),
    .X(_05999_));
 sg13g2_buf_2 fanout504 (.A(net507),
    .X(net504));
 sg13g2_mux4_1 _11999_ (.S0(net579),
    .A0(_05684_),
    .A1(_04278_),
    .A2(_05868_),
    .A3(_04177_),
    .S1(net589),
    .X(_06001_));
 sg13g2_buf_1 fanout503 (.A(net509),
    .X(net503));
 sg13g2_nor2_1 _12001_ (.A(net382),
    .B(_06001_),
    .Y(_06003_));
 sg13g2_a21o_1 _12002_ (.A2(_05999_),
    .A1(net382),
    .B1(_06003_),
    .X(_06004_));
 sg13g2_buf_1 fanout502 (.A(net503),
    .X(net502));
 sg13g2_nor2_1 _12004_ (.A(net364),
    .B(_06004_),
    .Y(_06006_));
 sg13g2_nor2_1 _12005_ (.A(net1253),
    .B(net823),
    .Y(_06007_));
 sg13g2_o21ai_1 _12006_ (.B1(_06007_),
    .Y(_06008_),
    .A1(_05998_),
    .A2(_06006_));
 sg13g2_a21o_1 _12007_ (.A2(net381),
    .A1(net628),
    .B1(net361),
    .X(_06009_));
 sg13g2_nor2_1 _12008_ (.A(_06003_),
    .B(_06009_),
    .Y(_06010_));
 sg13g2_o21ai_1 _12009_ (.B1(_05853_),
    .Y(_06011_),
    .A1(_05998_),
    .A2(_06010_));
 sg13g2_buf_2 fanout501 (.A(net503),
    .X(net501));
 sg13g2_a21oi_1 _12011_ (.A1(_06008_),
    .A2(_06011_),
    .Y(_06013_),
    .B1(net350));
 sg13g2_mux2_1 _12012_ (.A0(net391),
    .A1(_05842_),
    .S(net572),
    .X(_06014_));
 sg13g2_mux2_1 _12013_ (.A0(_05934_),
    .A1(_06014_),
    .S(net592),
    .X(_06015_));
 sg13g2_buf_2 fanout500 (.A(net503),
    .X(net500));
 sg13g2_nand2_1 _12015_ (.Y(_06017_),
    .A(_05818_),
    .B(_06015_));
 sg13g2_o21ai_1 _12016_ (.B1(net834),
    .Y(_06018_),
    .A1(_05790_),
    .A2(_06017_));
 sg13g2_a22oi_1 _12017_ (.Y(_06019_),
    .B1(_06013_),
    .B2(_06018_),
    .A2(_05993_),
    .A1(_05914_));
 sg13g2_and3_1 _12018_ (.X(_06020_),
    .A(net1240),
    .B(_03851_),
    .C(_03881_));
 sg13g2_buf_2 fanout499 (.A(net500),
    .X(net499));
 sg13g2_nor2_1 _12020_ (.A(net814),
    .B(net636),
    .Y(_06022_));
 sg13g2_buf_1 fanout498 (.A(_08312_),
    .X(net498));
 sg13g2_xnor2_1 _12022_ (.Y(_06024_),
    .A(_05458_),
    .B(_05498_));
 sg13g2_nand2_1 _12023_ (.Y(_06025_),
    .A(net596),
    .B(_05969_));
 sg13g2_o21ai_1 _12024_ (.B1(_06025_),
    .Y(_06026_),
    .A1(_05662_),
    .A2(_05971_));
 sg13g2_xnor2_1 _12025_ (.Y(_06027_),
    .A(_06024_),
    .B(_06026_));
 sg13g2_nor2_1 _12026_ (.A(net850),
    .B(_06024_),
    .Y(_06028_));
 sg13g2_buf_2 fanout497 (.A(net498),
    .X(net497));
 sg13g2_o21ai_1 _12028_ (.B1(net846),
    .Y(_06030_),
    .A1(net820),
    .A2(_05926_));
 sg13g2_nor2_1 _12029_ (.A(net845),
    .B(_05926_),
    .Y(_06031_));
 sg13g2_a21oi_1 _12030_ (.A1(_05458_),
    .A2(_06030_),
    .Y(_06032_),
    .B1(_06031_));
 sg13g2_o21ai_1 _12031_ (.B1(net839),
    .Y(_06033_),
    .A1(net565),
    .A2(_06032_));
 sg13g2_a22oi_1 _12032_ (.Y(_06034_),
    .B1(_06028_),
    .B2(_06033_),
    .A2(_06027_),
    .A1(net346));
 sg13g2_nor2_1 _12033_ (.A(_06019_),
    .B(_06034_),
    .Y(net91));
 sg13g2_a21oi_1 _12034_ (.A1(_05585_),
    .A2(_05598_),
    .Y(_06035_),
    .B1(_05662_));
 sg13g2_nand2_1 _12035_ (.Y(_06036_),
    .A(_05526_),
    .B(_05591_));
 sg13g2_nand2_1 _12036_ (.Y(_06037_),
    .A(net597),
    .B(_05458_));
 sg13g2_nand3b_1 _12037_ (.B(_06036_),
    .C(_06037_),
    .Y(_06038_),
    .A_N(_06035_));
 sg13g2_a21o_1 _12038_ (.A2(_06035_),
    .A1(_05573_),
    .B1(net912),
    .X(_06039_));
 sg13g2_a21oi_1 _12039_ (.A1(_06038_),
    .A2(_06039_),
    .Y(_06040_),
    .B1(_05436_));
 sg13g2_nor2_1 _12040_ (.A(_05566_),
    .B(_05665_),
    .Y(_06041_));
 sg13g2_nand2b_1 _12041_ (.Y(_06042_),
    .B(_06041_),
    .A_N(_06040_));
 sg13g2_nand2_1 _12042_ (.Y(_06043_),
    .A(net837),
    .B(net345));
 sg13g2_buf_2 fanout496 (.A(net497),
    .X(net496));
 sg13g2_buf_2 fanout495 (.A(net497),
    .X(net495));
 sg13g2_buf_1 fanout494 (.A(net495),
    .X(net494));
 sg13g2_o21ai_1 _12046_ (.B1(net814),
    .Y(_06047_),
    .A1(net611),
    .A2(_05290_));
 sg13g2_nand2_1 _12047_ (.Y(_06048_),
    .A(net850),
    .B(_05291_));
 sg13g2_a21oi_1 _12048_ (.A1(_06047_),
    .A2(_06048_),
    .Y(_06049_),
    .B1(net564));
 sg13g2_buf_2 fanout493 (.A(net497),
    .X(net493));
 sg13g2_mux4_1 _12050_ (.S0(net572),
    .A0(net611),
    .A1(net596),
    .A2(net391),
    .A3(_05842_),
    .S1(net644),
    .X(_06051_));
 sg13g2_nor2_1 _12051_ (.A(net373),
    .B(_05791_),
    .Y(_06052_));
 sg13g2_a21o_1 _12052_ (.A2(_06051_),
    .A1(net373),
    .B1(_06052_),
    .X(_06053_));
 sg13g2_buf_2 fanout492 (.A(net498),
    .X(net492));
 sg13g2_nor2_1 _12054_ (.A(net868),
    .B(_06053_),
    .Y(_06055_));
 sg13g2_a22oi_1 _12055_ (.Y(_06056_),
    .B1(_05761_),
    .B2(net375),
    .A2(_05756_),
    .A1(net594));
 sg13g2_a22oi_1 _12056_ (.Y(_06057_),
    .B1(_06056_),
    .B2(net824),
    .A2(_05772_),
    .A1(net375));
 sg13g2_nor3_1 _12057_ (.A(net399),
    .B(_06055_),
    .C(_06057_),
    .Y(_06058_));
 sg13g2_nor2_1 _12058_ (.A(net375),
    .B(_05727_),
    .Y(_06059_));
 sg13g2_a21oi_1 _12059_ (.A1(net375),
    .A2(_05750_),
    .Y(_06060_),
    .B1(_06059_));
 sg13g2_nor2_1 _12060_ (.A(net367),
    .B(net824),
    .Y(_06061_));
 sg13g2_nor2b_1 _12061_ (.A(_06060_),
    .B_N(_06061_),
    .Y(_06062_));
 sg13g2_nor3_1 _12062_ (.A(net608),
    .B(_06058_),
    .C(_06062_),
    .Y(_06063_));
 sg13g2_nor2_2 _12063_ (.A(net629),
    .B(_05956_),
    .Y(_06064_));
 sg13g2_buf_2 fanout491 (.A(net492),
    .X(net491));
 sg13g2_a21oi_1 _12065_ (.A1(net362),
    .A2(_05734_),
    .Y(_06066_),
    .B1(net373));
 sg13g2_nand2_1 _12066_ (.Y(_06067_),
    .A(net383),
    .B(_05734_));
 sg13g2_o21ai_1 _12067_ (.B1(_06067_),
    .Y(_06068_),
    .A1(net383),
    .A2(_05720_));
 sg13g2_nor2_1 _12068_ (.A(net395),
    .B(_06068_),
    .Y(_06069_));
 sg13g2_nor2_1 _12069_ (.A(net384),
    .B(net363),
    .Y(_06070_));
 sg13g2_nor2_1 _12070_ (.A(net823),
    .B(_05738_),
    .Y(_06071_));
 sg13g2_a21o_1 _12071_ (.A2(_06071_),
    .A1(_06070_),
    .B1(net348),
    .X(_06072_));
 sg13g2_a221oi_1 _12072_ (.B2(net870),
    .C1(_06072_),
    .B1(_06069_),
    .A1(_06064_),
    .Y(_06073_),
    .A2(_06066_));
 sg13g2_nor3_1 _12073_ (.A(net839),
    .B(_06063_),
    .C(_06073_),
    .Y(_06074_));
 sg13g2_a22oi_1 _12074_ (.Y(_06075_),
    .B1(_06049_),
    .B2(_06074_),
    .A2(_05436_),
    .A1(net820));
 sg13g2_o21ai_1 _12075_ (.B1(_06075_),
    .Y(net92),
    .A1(_06042_),
    .A2(_06043_));
 sg13g2_and3_2 _12076_ (.X(_06076_),
    .A(_05300_),
    .B(_05307_),
    .C(_05315_));
 sg13g2_buf_1 fanout490 (.A(net498),
    .X(net490));
 sg13g2_xnor2_1 _12078_ (.Y(_06078_),
    .A(_06076_),
    .B(_05322_));
 sg13g2_a21oi_1 _12079_ (.A1(net850),
    .A2(_06076_),
    .Y(_06079_),
    .B1(net814));
 sg13g2_nand2_1 _12080_ (.Y(_06080_),
    .A(net814),
    .B(_06076_));
 sg13g2_o21ai_1 _12081_ (.B1(_06080_),
    .Y(_06081_),
    .A1(_05322_),
    .A2(_06079_));
 sg13g2_a221oi_1 _12082_ (.B2(net636),
    .C1(net833),
    .B1(_06081_),
    .A1(net820),
    .Y(_06082_),
    .A2(_06078_));
 sg13g2_buf_2 fanout489 (.A(net498),
    .X(net489));
 sg13g2_nor3_1 _12084_ (.A(_05291_),
    .B(_05566_),
    .C(_05665_),
    .Y(_06084_));
 sg13g2_xnor2_1 _12085_ (.Y(_06085_),
    .A(_06078_),
    .B(_06084_));
 sg13g2_nand2_1 _12086_ (.Y(_06086_),
    .A(net346),
    .B(_06085_));
 sg13g2_mux4_1 _12087_ (.S0(net592),
    .A0(net611),
    .A1(_06076_),
    .A2(net596),
    .A3(net391),
    .S1(net573),
    .X(_06087_));
 sg13g2_mux2_1 _12088_ (.A0(_05822_),
    .A1(_06087_),
    .S(net375),
    .X(_06088_));
 sg13g2_nor2_1 _12089_ (.A(net375),
    .B(_05834_),
    .Y(_06089_));
 sg13g2_a22oi_1 _12090_ (.Y(_06090_),
    .B1(_06089_),
    .B2(net824),
    .A2(_05847_),
    .A1(net376));
 sg13g2_a21oi_1 _12091_ (.A1(net824),
    .A2(_06088_),
    .Y(_06091_),
    .B1(_06090_));
 sg13g2_nor2_1 _12092_ (.A(net387),
    .B(_05838_),
    .Y(_06092_));
 sg13g2_a21oi_1 _12093_ (.A1(net387),
    .A2(_05857_),
    .Y(_06093_),
    .B1(_06092_));
 sg13g2_nand2_1 _12094_ (.Y(_06094_),
    .A(_06061_),
    .B(_06093_));
 sg13g2_o21ai_1 _12095_ (.B1(_06094_),
    .Y(_06095_),
    .A1(net399),
    .A2(_06091_));
 sg13g2_nand2_1 _12096_ (.Y(_06096_),
    .A(net369),
    .B(net392));
 sg13g2_nor2_1 _12097_ (.A(net381),
    .B(_05860_),
    .Y(_06097_));
 sg13g2_a21oi_1 _12098_ (.A1(net381),
    .A2(_05864_),
    .Y(_06098_),
    .B1(_06097_));
 sg13g2_nand2_1 _12099_ (.Y(_06099_),
    .A(net361),
    .B(_06098_));
 sg13g2_o21ai_1 _12100_ (.B1(_06099_),
    .Y(_06100_),
    .A1(_06096_),
    .A2(_05884_));
 sg13g2_nor3_1 _12101_ (.A(net381),
    .B(_05867_),
    .C(_05871_),
    .Y(_06101_));
 sg13g2_nor2_1 _12102_ (.A(_06009_),
    .B(_06101_),
    .Y(_06102_));
 sg13g2_a21oi_1 _12103_ (.A1(net361),
    .A2(_06098_),
    .Y(_06103_),
    .B1(_06102_));
 sg13g2_nand2_1 _12104_ (.Y(_06104_),
    .A(net1253),
    .B(_06103_));
 sg13g2_o21ai_1 _12105_ (.B1(_06104_),
    .Y(_06105_),
    .A1(net1253),
    .A2(_06100_));
 sg13g2_nor3_1 _12106_ (.A(net351),
    .B(net825),
    .C(_06105_),
    .Y(_06106_));
 sg13g2_buf_2 fanout488 (.A(net490),
    .X(net488));
 sg13g2_a22oi_1 _12108_ (.Y(_06108_),
    .B1(_06106_),
    .B2(net838),
    .A2(_06095_),
    .A1(net351));
 sg13g2_a21oi_1 _12109_ (.A1(_06082_),
    .A2(_06086_),
    .Y(net93),
    .B1(_06108_));
 sg13g2_nor2_1 _12110_ (.A(net387),
    .B(_05924_),
    .Y(_06109_));
 sg13g2_a21oi_1 _12111_ (.A1(net387),
    .A2(_05948_),
    .Y(_06110_),
    .B1(_06109_));
 sg13g2_buf_2 fanout487 (.A(_08389_),
    .X(net487));
 sg13g2_mux4_1 _12113_ (.S0(net583),
    .A0(net611),
    .A1(net599),
    .A2(net391),
    .A3(_06076_),
    .S1(net644),
    .X(_06112_));
 sg13g2_mux2_1 _12114_ (.A0(_05936_),
    .A1(_06112_),
    .S(net375),
    .X(_06113_));
 sg13g2_nor2_1 _12115_ (.A(net868),
    .B(_06113_),
    .Y(_06114_));
 sg13g2_nor2_1 _12116_ (.A(net389),
    .B(_05930_),
    .Y(_06115_));
 sg13g2_a22oi_1 _12117_ (.Y(_06116_),
    .B1(_06115_),
    .B2(net824),
    .A2(_05920_),
    .A1(net388));
 sg13g2_nor3_1 _12118_ (.A(net399),
    .B(_06114_),
    .C(_06116_),
    .Y(_06117_));
 sg13g2_a22oi_1 _12119_ (.Y(_06118_),
    .B1(_06117_),
    .B2(net608),
    .A2(_06110_),
    .A1(_06061_));
 sg13g2_nand2_1 _12120_ (.Y(_06119_),
    .A(net370),
    .B(net580));
 sg13g2_nor2_1 _12121_ (.A(net627),
    .B(net361),
    .Y(_06120_));
 sg13g2_nor2_1 _12122_ (.A(net570),
    .B(_05939_),
    .Y(_06121_));
 sg13g2_a21oi_1 _12123_ (.A1(net392),
    .A2(_06121_),
    .Y(_06122_),
    .B1(_05959_));
 sg13g2_nor2_1 _12124_ (.A(net374),
    .B(net396),
    .Y(_06123_));
 sg13g2_nand2_1 _12125_ (.Y(_06124_),
    .A(_06123_),
    .B(_05944_));
 sg13g2_o21ai_1 _12126_ (.B1(_06124_),
    .Y(_06125_),
    .A1(net380),
    .A2(_06122_));
 sg13g2_a21o_1 _12127_ (.A2(_06120_),
    .A1(_06119_),
    .B1(_06125_),
    .X(_06126_));
 sg13g2_and2_1 _12128_ (.A(_06007_),
    .B(_06125_),
    .X(_06127_));
 sg13g2_a22oi_1 _12129_ (.Y(_06128_),
    .B1(_06127_),
    .B2(net349),
    .A2(_06126_),
    .A1(_05853_));
 sg13g2_or2_1 _12130_ (.X(_06129_),
    .B(_06128_),
    .A(_06118_));
 sg13g2_nor2_1 _12131_ (.A(_05291_),
    .B(_06076_),
    .Y(_06130_));
 sg13g2_and2_1 _12132_ (.A(net604),
    .B(_05322_),
    .X(_06131_));
 sg13g2_a221oi_1 _12133_ (.B2(_06041_),
    .C1(_06131_),
    .B1(_06130_),
    .A1(_05322_),
    .Y(_06132_),
    .A2(_06084_));
 sg13g2_xnor2_1 _12134_ (.Y(_06133_),
    .A(_05429_),
    .B(_06132_));
 sg13g2_o21ai_1 _12135_ (.B1(net845),
    .Y(_06134_),
    .A1(net820),
    .A2(net602));
 sg13g2_buf_2 fanout486 (.A(net487),
    .X(net486));
 sg13g2_nor2_1 _12137_ (.A(net845),
    .B(_05411_),
    .Y(_06136_));
 sg13g2_a21oi_1 _12138_ (.A1(_05426_),
    .A2(_06134_),
    .Y(_06137_),
    .B1(_06136_));
 sg13g2_o21ai_1 _12139_ (.B1(net839),
    .Y(_06138_),
    .A1(net564),
    .A2(_06137_));
 sg13g2_nor2_1 _12140_ (.A(net850),
    .B(_05429_),
    .Y(_06139_));
 sg13g2_a22oi_1 _12141_ (.Y(_06140_),
    .B1(_06138_),
    .B2(_06139_),
    .A2(_06133_),
    .A1(net346));
 sg13g2_a21oi_1 _12142_ (.A1(net834),
    .A2(_06129_),
    .Y(net94),
    .B1(_06140_));
 sg13g2_nor2_1 _12143_ (.A(net833),
    .B(net357),
    .Y(_06141_));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_nor2b_1 _12145_ (.A(_05413_),
    .B_N(_05423_),
    .Y(_06143_));
 sg13g2_nor2_1 _12146_ (.A(_05426_),
    .B(net599),
    .Y(_06144_));
 sg13g2_nor2_1 _12147_ (.A(_06144_),
    .B(_05423_),
    .Y(_06145_));
 sg13g2_mux2_1 _12148_ (.A0(_06143_),
    .A1(_06145_),
    .S(_06132_),
    .X(_06146_));
 sg13g2_mux2_1 _12149_ (.A0(_05413_),
    .A1(_06144_),
    .S(_05423_),
    .X(_06147_));
 sg13g2_nor2_1 _12150_ (.A(_05333_),
    .B(_05362_),
    .Y(_06148_));
 sg13g2_nand3_1 _12151_ (.B(_05333_),
    .C(_05362_),
    .A(net850),
    .Y(_06149_));
 sg13g2_o21ai_1 _12152_ (.B1(_06149_),
    .Y(_06150_),
    .A1(net845),
    .A2(_06148_));
 sg13g2_and2_1 _12153_ (.A(net636),
    .B(_06150_),
    .X(_06151_));
 sg13g2_a221oi_1 _12154_ (.B2(_06147_),
    .C1(_06151_),
    .B1(net346),
    .A1(net820),
    .Y(_06152_),
    .A2(_05423_));
 sg13g2_mux2_1 _12155_ (.A0(_05980_),
    .A1(_05986_),
    .S(net366),
    .X(_06153_));
 sg13g2_and2_1 _12156_ (.A(net399),
    .B(_05994_),
    .X(_06154_));
 sg13g2_a22oi_1 _12157_ (.Y(_06155_),
    .B1(_06154_),
    .B2(net376),
    .A2(_05981_),
    .A1(net367));
 sg13g2_a22oi_1 _12158_ (.Y(_06156_),
    .B1(_06155_),
    .B2(net824),
    .A2(_06153_),
    .A1(net376));
 sg13g2_mux4_1 _12159_ (.S0(net591),
    .A0(_05434_),
    .A1(net603),
    .A2(net602),
    .A3(net600),
    .S1(net582),
    .X(_06157_));
 sg13g2_nor2_1 _12160_ (.A(net384),
    .B(_06157_),
    .Y(_06158_));
 sg13g2_a21oi_1 _12161_ (.A1(net384),
    .A2(_06015_),
    .Y(_06159_),
    .B1(_06158_));
 sg13g2_nor3_1 _12162_ (.A(net396),
    .B(net868),
    .C(_06159_),
    .Y(_06160_));
 sg13g2_or2_1 _12163_ (.X(_06161_),
    .B(_06160_),
    .A(_06156_));
 sg13g2_nand2_1 _12164_ (.Y(_06162_),
    .A(net371),
    .B(_05995_));
 sg13g2_o21ai_1 _12165_ (.B1(_06162_),
    .Y(_06163_),
    .A1(net370),
    .A2(_06001_));
 sg13g2_buf_2 fanout484 (.A(net486),
    .X(net484));
 sg13g2_nor2_1 _12167_ (.A(_04391_),
    .B(net628),
    .Y(_06165_));
 sg13g2_nor3_1 _12168_ (.A(net1253),
    .B(net385),
    .C(_05999_),
    .Y(_06166_));
 sg13g2_nor3_1 _12169_ (.A(net364),
    .B(_06165_),
    .C(_06166_),
    .Y(_06167_));
 sg13g2_a22oi_1 _12170_ (.Y(_06168_),
    .B1(_06167_),
    .B2(net826),
    .A2(_06163_),
    .A1(net364));
 sg13g2_and2_1 _12171_ (.A(net609),
    .B(_06168_),
    .X(_06169_));
 sg13g2_a22oi_1 _12172_ (.Y(_06170_),
    .B1(_06169_),
    .B2(net838),
    .A2(_06161_),
    .A1(net351));
 sg13g2_a21oi_1 _12173_ (.A1(net839),
    .A2(_06152_),
    .Y(_06171_),
    .B1(_06170_));
 sg13g2_a21o_1 _12174_ (.A2(_06146_),
    .A1(_06141_),
    .B1(_06171_),
    .X(net95));
 sg13g2_o21ai_1 _12175_ (.B1(_05419_),
    .Y(_06172_),
    .A1(_06041_),
    .A2(_05431_));
 sg13g2_buf_2 fanout483 (.A(net484),
    .X(net483));
 sg13g2_nor3_1 _12177_ (.A(net814),
    .B(net821),
    .C(net614),
    .Y(_06174_));
 sg13g2_nand3_1 _12178_ (.B(_06172_),
    .C(_06174_),
    .A(_05239_),
    .Y(_06175_));
 sg13g2_nor4_1 _12179_ (.A(net814),
    .B(net636),
    .C(net614),
    .D(_05239_),
    .Y(_06176_));
 sg13g2_nand2b_1 _12180_ (.Y(_06177_),
    .B(_06176_),
    .A_N(_06172_));
 sg13g2_nor4_1 _12181_ (.A(net564),
    .B(net614),
    .C(_05030_),
    .D(_05034_),
    .Y(_06178_));
 sg13g2_nor3_1 _12182_ (.A(net851),
    .B(net614),
    .C(_05239_),
    .Y(_06179_));
 sg13g2_nor3_1 _12183_ (.A(net846),
    .B(net564),
    .C(net614),
    .Y(_06180_));
 sg13g2_a22oi_1 _12184_ (.Y(_06181_),
    .B1(_06179_),
    .B2(_06180_),
    .A2(_06178_),
    .A1(net851));
 sg13g2_nand3_1 _12185_ (.B(_06177_),
    .C(_06181_),
    .A(_06175_),
    .Y(_06182_));
 sg13g2_nor4_1 _12186_ (.A(net851),
    .B(_05237_),
    .C(_05030_),
    .D(_05034_),
    .Y(_06183_));
 sg13g2_xnor2_1 _12187_ (.Y(_06184_),
    .A(_05239_),
    .B(_06172_));
 sg13g2_nor3_1 _12188_ (.A(_05237_),
    .B(net357),
    .C(_06184_),
    .Y(_06185_));
 sg13g2_nor2_1 _12189_ (.A(net846),
    .B(net564),
    .Y(_06186_));
 sg13g2_and2_1 _12190_ (.A(_05239_),
    .B(_06186_),
    .X(_06187_));
 sg13g2_nor4_1 _12191_ (.A(_06182_),
    .B(_06183_),
    .C(_06185_),
    .D(_06187_),
    .Y(_06188_));
 sg13g2_nor2_1 _12192_ (.A(net826),
    .B(_05739_),
    .Y(_06189_));
 sg13g2_buf_1 fanout482 (.A(net487),
    .X(net482));
 sg13g2_mux2_1 _12194_ (.A0(_06064_),
    .A1(_06189_),
    .S(net365),
    .X(_06191_));
 sg13g2_buf_2 fanout481 (.A(net482),
    .X(net481));
 sg13g2_mux4_1 _12196_ (.S0(net572),
    .A0(net613),
    .A1(net602),
    .A2(net600),
    .A3(net603),
    .S1(net643),
    .X(_06193_));
 sg13g2_nand2_1 _12197_ (.Y(_06194_),
    .A(net384),
    .B(_06051_));
 sg13g2_o21ai_1 _12198_ (.B1(_06194_),
    .Y(_06195_),
    .A1(net383),
    .A2(_06193_));
 sg13g2_nor2_1 _12199_ (.A(_06096_),
    .B(_05791_),
    .Y(_06196_));
 sg13g2_a21oi_1 _12200_ (.A1(net362),
    .A2(_06195_),
    .Y(_06197_),
    .B1(_06196_));
 sg13g2_nand2_1 _12201_ (.Y(_06198_),
    .A(net367),
    .B(_05763_));
 sg13g2_nand2_1 _12202_ (.Y(_06199_),
    .A(net395),
    .B(_05729_));
 sg13g2_a21oi_1 _12203_ (.A1(_06198_),
    .A2(_06199_),
    .Y(_06200_),
    .B1(_05912_));
 sg13g2_a22oi_1 _12204_ (.Y(_06201_),
    .B1(_06200_),
    .B2(net836),
    .A2(_06197_),
    .A1(net358));
 sg13g2_o21ai_1 _12205_ (.B1(_06201_),
    .Y(_06202_),
    .A1(net350),
    .A2(_06191_));
 sg13g2_o21ai_1 _12206_ (.B1(_06202_),
    .Y(net96),
    .A1(net834),
    .A2(_06188_));
 sg13g2_mux4_1 _12207_ (.S0(net591),
    .A0(net613),
    .A1(net566),
    .A2(net602),
    .A3(net600),
    .S1(net572),
    .X(_06203_));
 sg13g2_nor2_1 _12208_ (.A(net399),
    .B(_06203_),
    .Y(_06204_));
 sg13g2_a21oi_1 _12209_ (.A1(net399),
    .A2(_05822_),
    .Y(_06205_),
    .B1(_06204_));
 sg13g2_nand2_1 _12210_ (.Y(_06206_),
    .A(_06123_),
    .B(_06087_));
 sg13g2_o21ai_1 _12211_ (.B1(_06206_),
    .Y(_06207_),
    .A1(net387),
    .A2(_06205_));
 sg13g2_nor2_1 _12212_ (.A(net400),
    .B(_05840_),
    .Y(_06208_));
 sg13g2_a22oi_1 _12213_ (.Y(_06209_),
    .B1(_06208_),
    .B2(net609),
    .A2(_05862_),
    .A1(net397));
 sg13g2_nor2_1 _12214_ (.A(net1253),
    .B(net397),
    .Y(_06210_));
 sg13g2_a21o_1 _12215_ (.A2(_05871_),
    .A1(net361),
    .B1(_05867_),
    .X(_06211_));
 sg13g2_nor2_1 _12216_ (.A(net342),
    .B(_05864_),
    .Y(_06212_));
 sg13g2_a22oi_1 _12217_ (.Y(_06213_),
    .B1(_06212_),
    .B2(_06120_),
    .A2(_06211_),
    .A1(net381));
 sg13g2_nor2_1 _12218_ (.A(_04391_),
    .B(_06213_),
    .Y(_06214_));
 sg13g2_a22oi_1 _12219_ (.Y(_06215_),
    .B1(_06214_),
    .B2(net350),
    .A2(_06210_),
    .A1(_05886_));
 sg13g2_nor3_1 _12220_ (.A(net825),
    .B(_06209_),
    .C(_06215_),
    .Y(_06216_));
 sg13g2_a22oi_1 _12221_ (.Y(_06217_),
    .B1(_06216_),
    .B2(net838),
    .A2(_06207_),
    .A1(net358));
 sg13g2_xnor2_1 _12222_ (.Y(_06218_),
    .A(_04990_),
    .B(net566));
 sg13g2_o21ai_1 _12223_ (.B1(net846),
    .Y(_06219_),
    .A1(net821),
    .A2(net567));
 sg13g2_nand2_1 _12224_ (.Y(_06220_),
    .A(_04990_),
    .B(_06219_));
 sg13g2_o21ai_1 _12225_ (.B1(_06220_),
    .Y(_06221_),
    .A1(net846),
    .A2(net567));
 sg13g2_a221oi_1 _12226_ (.B2(net637),
    .C1(net833),
    .B1(_06221_),
    .A1(net821),
    .Y(_06222_),
    .A2(_06218_));
 sg13g2_nor2_1 _12227_ (.A(_05036_),
    .B(_05236_),
    .Y(_06223_));
 sg13g2_nor2_1 _12228_ (.A(_05237_),
    .B(_05239_),
    .Y(_06224_));
 sg13g2_nor2_1 _12229_ (.A(_06218_),
    .B(_06224_),
    .Y(_06225_));
 sg13g2_mux2_1 _12230_ (.A0(_06223_),
    .A1(_06225_),
    .S(_06172_),
    .X(_06226_));
 sg13g2_mux2_1 _12231_ (.A0(_05036_),
    .A1(_06224_),
    .S(_06218_),
    .X(_06227_));
 sg13g2_o21ai_1 _12232_ (.B1(net346),
    .Y(_06228_),
    .A1(_06226_),
    .A2(_06227_));
 sg13g2_and2_1 _12233_ (.A(_06222_),
    .B(_06228_),
    .X(_06229_));
 sg13g2_nor2_1 _12234_ (.A(_06217_),
    .B(_06229_),
    .Y(net97));
 sg13g2_nor2_1 _12235_ (.A(_05236_),
    .B(_05241_),
    .Y(_06230_));
 sg13g2_and2_1 _12236_ (.A(_06230_),
    .B(_06172_),
    .X(_06231_));
 sg13g2_nand2_1 _12237_ (.Y(_06232_),
    .A(_04990_),
    .B(_05036_));
 sg13g2_o21ai_1 _12238_ (.B1(_05120_),
    .Y(_06233_),
    .A1(_04990_),
    .A2(_05036_));
 sg13g2_nand2_1 _12239_ (.Y(_06234_),
    .A(_06232_),
    .B(_06233_));
 sg13g2_a21oi_1 _12240_ (.A1(_06230_),
    .A2(_06172_),
    .Y(_06235_),
    .B1(_06234_));
 sg13g2_xnor2_1 _12241_ (.Y(_06236_),
    .A(_05829_),
    .B(_04985_));
 sg13g2_mux2_1 _12242_ (.A0(_06231_),
    .A1(_06235_),
    .S(_06236_),
    .X(_06237_));
 sg13g2_nand2_1 _12243_ (.Y(_06238_),
    .A(net354),
    .B(_04986_));
 sg13g2_nand2_1 _12244_ (.Y(_06239_),
    .A(net814),
    .B(_06238_));
 sg13g2_o21ai_1 _12245_ (.B1(_06239_),
    .Y(_06240_),
    .A1(net820),
    .A2(_05089_));
 sg13g2_a21oi_1 _12246_ (.A1(net339),
    .A2(_06234_),
    .Y(_06241_),
    .B1(_06236_));
 sg13g2_a21oi_1 _12247_ (.A1(net851),
    .A2(_06236_),
    .Y(_06242_),
    .B1(_06241_));
 sg13g2_a21oi_1 _12248_ (.A1(net637),
    .A2(_06240_),
    .Y(_06243_),
    .B1(_06242_));
 sg13g2_o21ai_1 _12249_ (.B1(_05866_),
    .Y(_06244_),
    .A1(net394),
    .A2(_05940_));
 sg13g2_a221oi_1 _12250_ (.B2(net381),
    .C1(_06120_),
    .B1(_06244_),
    .A1(net341),
    .Y(_06245_),
    .A2(_05944_));
 sg13g2_nand2_1 _12251_ (.Y(_06246_),
    .A(_05947_),
    .B(_06210_));
 sg13g2_o21ai_1 _12252_ (.B1(_06246_),
    .Y(_06247_),
    .A1(_04391_),
    .A2(_06245_));
 sg13g2_and2_1 _12253_ (.A(net869),
    .B(_06247_),
    .X(_06248_));
 sg13g2_mux4_1 _12254_ (.S0(net582),
    .A0(net613),
    .A1(net354),
    .A2(net600),
    .A3(net566),
    .S1(net643),
    .X(_06249_));
 sg13g2_nor2_1 _12255_ (.A(net367),
    .B(_05936_),
    .Y(_06250_));
 sg13g2_a22oi_1 _12256_ (.Y(_06251_),
    .B1(_06250_),
    .B2(net387),
    .A2(_06249_),
    .A1(net367));
 sg13g2_a21oi_1 _12257_ (.A1(_06123_),
    .A2(_06112_),
    .Y(_06252_),
    .B1(_06251_));
 sg13g2_a21oi_1 _12258_ (.A1(net825),
    .A2(_06252_),
    .Y(_06253_),
    .B1(net609));
 sg13g2_nor2_1 _12259_ (.A(net366),
    .B(_05952_),
    .Y(_06254_));
 sg13g2_a22oi_1 _12260_ (.Y(_06255_),
    .B1(_06254_),
    .B2(_05912_),
    .A2(_05925_),
    .A1(net366));
 sg13g2_nor2_1 _12261_ (.A(net838),
    .B(_06255_),
    .Y(_06256_));
 sg13g2_o21ai_1 _12262_ (.B1(_06256_),
    .Y(_06257_),
    .A1(_06248_),
    .A2(_06253_));
 sg13g2_nand2_1 _12263_ (.Y(_06258_),
    .A(_06243_),
    .B(_06257_));
 sg13g2_a21o_1 _12264_ (.A2(_06237_),
    .A1(net339),
    .B1(_06258_),
    .X(net67));
 sg13g2_nand2_1 _12265_ (.Y(_06259_),
    .A(_05234_),
    .B(_06238_));
 sg13g2_nand2b_1 _12266_ (.Y(_06260_),
    .B(_05089_),
    .A_N(_05234_));
 sg13g2_mux2_1 _12267_ (.A0(_06259_),
    .A1(_06260_),
    .S(_06235_),
    .X(_06261_));
 sg13g2_mux4_1 _12268_ (.S0(net643),
    .A0(_05917_),
    .A1(net354),
    .A2(net566),
    .A3(net613),
    .S1(net573),
    .X(_06262_));
 sg13g2_mux2_1 _12269_ (.A0(_06157_),
    .A1(_06262_),
    .S(net372),
    .X(_06263_));
 sg13g2_nor2_1 _12270_ (.A(net396),
    .B(_06263_),
    .Y(_06264_));
 sg13g2_a21oi_1 _12271_ (.A1(_06070_),
    .A2(_06015_),
    .Y(_06265_),
    .B1(_06264_));
 sg13g2_nor2_1 _12272_ (.A(net366),
    .B(_05997_),
    .Y(_06266_));
 sg13g2_a22oi_1 _12273_ (.Y(_06267_),
    .B1(_06266_),
    .B2(_05912_),
    .A2(_05983_),
    .A1(net366));
 sg13g2_a21oi_1 _12274_ (.A1(net358),
    .A2(_06265_),
    .Y(_06268_),
    .B1(_06267_));
 sg13g2_nor2_1 _12275_ (.A(_05793_),
    .B(_06001_),
    .Y(_06269_));
 sg13g2_a22oi_1 _12276_ (.Y(_06270_),
    .B1(_05956_),
    .B2(_06269_),
    .A2(_05793_),
    .A1(net628));
 sg13g2_nor3_1 _12277_ (.A(net394),
    .B(_05888_),
    .C(_06004_),
    .Y(_06271_));
 sg13g2_nor3_1 _12278_ (.A(net349),
    .B(_06270_),
    .C(_06271_),
    .Y(_06272_));
 sg13g2_nor2_1 _12279_ (.A(net839),
    .B(_06272_),
    .Y(_06273_));
 sg13g2_mux2_1 _12280_ (.A0(_06238_),
    .A1(_05089_),
    .S(_05234_),
    .X(_06274_));
 sg13g2_nor2_1 _12281_ (.A(_06043_),
    .B(_06274_),
    .Y(_06275_));
 sg13g2_nand2_1 _12282_ (.Y(_06276_),
    .A(net851),
    .B(_05174_));
 sg13g2_o21ai_1 _12283_ (.B1(_06276_),
    .Y(_06277_),
    .A1(net846),
    .A2(_05172_));
 sg13g2_nand2_1 _12284_ (.Y(_06278_),
    .A(net636),
    .B(_06277_));
 sg13g2_o21ai_1 _12285_ (.B1(_06278_),
    .Y(_06279_),
    .A1(net850),
    .A2(_05234_));
 sg13g2_a22oi_1 _12286_ (.Y(_06280_),
    .B1(_06275_),
    .B2(_06279_),
    .A2(_06273_),
    .A1(_06268_));
 sg13g2_o21ai_1 _12287_ (.B1(_06280_),
    .Y(net68),
    .A1(net340),
    .A2(_06261_));
 sg13g2_a21oi_1 _12288_ (.A1(net402),
    .A2(net573),
    .Y(_06281_),
    .B1(_05746_));
 sg13g2_a22oi_1 _12289_ (.Y(_06282_),
    .B1(_05984_),
    .B2(net594),
    .A2(net584),
    .A1(net401));
 sg13g2_a21oi_1 _12290_ (.A1(net593),
    .A2(_06281_),
    .Y(_06283_),
    .B1(_06282_));
 sg13g2_nor2_1 _12291_ (.A(net373),
    .B(_06193_),
    .Y(_06284_));
 sg13g2_a21oi_1 _12292_ (.A1(net373),
    .A2(_06283_),
    .Y(_06285_),
    .B1(_06284_));
 sg13g2_nor2_1 _12293_ (.A(net362),
    .B(_06053_),
    .Y(_06286_));
 sg13g2_a21oi_1 _12294_ (.A1(net362),
    .A2(_06285_),
    .Y(_06287_),
    .B1(_06286_));
 sg13g2_o21ai_1 _12295_ (.B1(net348),
    .Y(_06288_),
    .A1(net870),
    .A2(_06287_));
 sg13g2_a21o_1 _12296_ (.A2(net610),
    .A1(net628),
    .B1(_05956_),
    .X(_06289_));
 sg13g2_buf_2 fanout480 (.A(net482),
    .X(net480));
 sg13g2_nor3_1 _12298_ (.A(net348),
    .B(net341),
    .C(net343),
    .Y(_06291_));
 sg13g2_a21oi_1 _12299_ (.A1(net341),
    .A2(_06071_),
    .Y(_06292_),
    .B1(_06291_));
 sg13g2_nand2_1 _12300_ (.Y(_06293_),
    .A(_06288_),
    .B(_06292_));
 sg13g2_mux2_1 _12301_ (.A0(_06060_),
    .A1(_06068_),
    .S(net399),
    .X(_06294_));
 sg13g2_nand2_1 _12302_ (.Y(_06295_),
    .A(_05914_),
    .B(_06294_));
 sg13g2_a21oi_1 _12303_ (.A1(_06293_),
    .A2(_06295_),
    .Y(_06296_),
    .B1(net838));
 sg13g2_xnor2_1 _12304_ (.Y(_06297_),
    .A(net875),
    .B(_04976_));
 sg13g2_nand4_1 _12305_ (.B(net851),
    .C(net615),
    .A(net846),
    .Y(_06298_),
    .D(_06297_));
 sg13g2_or2_1 _12306_ (.X(_06299_),
    .B(net615),
    .A(net636));
 sg13g2_nand3b_1 _12307_ (.B(net847),
    .C(net403),
    .Y(_06300_),
    .A_N(_06299_));
 sg13g2_and3_1 _12308_ (.X(_06301_),
    .A(_05242_),
    .B(_05423_),
    .C(_05430_));
 sg13g2_o21ai_1 _12309_ (.B1(_06301_),
    .Y(_06302_),
    .A1(_05566_),
    .A2(_05665_));
 sg13g2_buf_2 fanout479 (.A(net480),
    .X(net479));
 sg13g2_a21oi_2 _12311_ (.B1(_05175_),
    .Y(_06304_),
    .A2(_05433_),
    .A1(_05242_));
 sg13g2_and2_1 _12312_ (.A(_06302_),
    .B(_06304_),
    .X(_06305_));
 sg13g2_a21oi_1 _12313_ (.A1(_06298_),
    .A2(_06300_),
    .Y(_06306_),
    .B1(_06305_));
 sg13g2_nand2_1 _12314_ (.Y(_06307_),
    .A(_06302_),
    .B(_06304_));
 sg13g2_nor4_1 _12315_ (.A(_06020_),
    .B(net403),
    .C(_06307_),
    .D(_06299_),
    .Y(_06308_));
 sg13g2_nand4_1 _12316_ (.B(net564),
    .C(net615),
    .A(net847),
    .Y(_06309_),
    .D(_04977_));
 sg13g2_and2_1 _12317_ (.A(net637),
    .B(net616),
    .X(_06310_));
 sg13g2_nand2b_1 _12318_ (.Y(_06311_),
    .B(net821),
    .A_N(net615));
 sg13g2_nand2_1 _12319_ (.Y(_06312_),
    .A(net851),
    .B(_06310_));
 sg13g2_a21oi_1 _12320_ (.A1(_06311_),
    .A2(_06312_),
    .Y(_06313_),
    .B1(net403));
 sg13g2_nand2_1 _12321_ (.Y(_06314_),
    .A(_06297_),
    .B(_06186_));
 sg13g2_nand3_1 _12322_ (.B(net615),
    .C(net403),
    .A(net821),
    .Y(_06315_));
 sg13g2_nand2_1 _12323_ (.Y(_06316_),
    .A(_06314_),
    .B(_06315_));
 sg13g2_a22oi_1 _12324_ (.Y(_06317_),
    .B1(_06313_),
    .B2(_06316_),
    .A2(_06310_),
    .A1(net814));
 sg13g2_o21ai_1 _12325_ (.B1(_06317_),
    .Y(_06318_),
    .A1(_06307_),
    .A2(_06309_));
 sg13g2_nor4_1 _12326_ (.A(net833),
    .B(_06306_),
    .C(_06308_),
    .D(_06318_),
    .Y(_06319_));
 sg13g2_nor2_1 _12327_ (.A(_06296_),
    .B(_06319_),
    .Y(net69));
 sg13g2_nand3_1 _12328_ (.B(_06302_),
    .C(_06304_),
    .A(net403),
    .Y(_06320_));
 sg13g2_a21oi_1 _12329_ (.A1(_06302_),
    .A2(_06304_),
    .Y(_06321_),
    .B1(net403));
 sg13g2_a21o_1 _12330_ (.A2(_06320_),
    .A1(net615),
    .B1(_06321_),
    .X(_06322_));
 sg13g2_xnor2_1 _12331_ (.Y(_06323_),
    .A(_04934_),
    .B(_06322_));
 sg13g2_and2_1 _12332_ (.A(_05185_),
    .B(_04933_),
    .X(_06324_));
 sg13g2_buf_2 fanout478 (.A(net480),
    .X(net478));
 sg13g2_nand2_1 _12334_ (.Y(_06326_),
    .A(net852),
    .B(_05192_));
 sg13g2_o21ai_1 _12335_ (.B1(_06326_),
    .Y(_06327_),
    .A1(net847),
    .A2(_06324_));
 sg13g2_mux2_1 _12336_ (.A0(_05185_),
    .A1(_05917_),
    .S(net573),
    .X(_06328_));
 sg13g2_a22oi_1 _12337_ (.Y(_06329_),
    .B1(_05746_),
    .B2(net593),
    .A2(net573),
    .A1(net402));
 sg13g2_a21oi_1 _12338_ (.A1(net593),
    .A2(_06328_),
    .Y(_06330_),
    .B1(_06329_));
 sg13g2_nor2_1 _12339_ (.A(net372),
    .B(_06203_),
    .Y(_06331_));
 sg13g2_a21oi_1 _12340_ (.A1(net372),
    .A2(_06330_),
    .Y(_06332_),
    .B1(_06331_));
 sg13g2_nor2_1 _12341_ (.A(net395),
    .B(_06332_),
    .Y(_06333_));
 sg13g2_a21oi_1 _12342_ (.A1(net395),
    .A2(_06088_),
    .Y(_06334_),
    .B1(_06333_));
 sg13g2_a21oi_1 _12343_ (.A1(net580),
    .A2(net341),
    .Y(_06335_),
    .B1(net627));
 sg13g2_a21oi_1 _12344_ (.A1(net341),
    .A2(_05871_),
    .Y(_06336_),
    .B1(_06335_));
 sg13g2_nor3_1 _12345_ (.A(net342),
    .B(_05888_),
    .C(_05884_),
    .Y(_06337_));
 sg13g2_nor2_1 _12346_ (.A(net349),
    .B(_06337_),
    .Y(_06338_));
 sg13g2_o21ai_1 _12347_ (.B1(_06338_),
    .Y(_06339_),
    .A1(_05956_),
    .A2(_06336_));
 sg13g2_nand2_1 _12348_ (.Y(_06340_),
    .A(net831),
    .B(_06339_));
 sg13g2_and2_1 _12349_ (.A(net366),
    .B(_06093_),
    .X(_06341_));
 sg13g2_a22oi_1 _12350_ (.Y(_06342_),
    .B1(_06341_),
    .B2(_05912_),
    .A2(_06098_),
    .A1(net398));
 sg13g2_a22oi_1 _12351_ (.Y(_06343_),
    .B1(_06340_),
    .B2(_06342_),
    .A2(_06334_),
    .A1(net358));
 sg13g2_a221oi_1 _12352_ (.B2(net637),
    .C1(_06343_),
    .B1(_06327_),
    .A1(net821),
    .Y(_06344_),
    .A2(_04934_));
 sg13g2_o21ai_1 _12353_ (.B1(_06344_),
    .Y(net70),
    .A1(net340),
    .A2(_06323_));
 sg13g2_nor2b_1 _12354_ (.A(_06324_),
    .B_N(net615),
    .Y(_06345_));
 sg13g2_a22oi_1 _12355_ (.Y(_06346_),
    .B1(net403),
    .B2(_06324_),
    .A2(_06304_),
    .A1(_06302_));
 sg13g2_a22oi_1 _12356_ (.Y(_06347_),
    .B1(_06346_),
    .B2(_05192_),
    .A2(_06345_),
    .A1(_06320_));
 sg13g2_xnor2_1 _12357_ (.Y(_06348_),
    .A(_04885_),
    .B(_06347_));
 sg13g2_nor2_1 _12358_ (.A(net360),
    .B(_06113_),
    .Y(_06349_));
 sg13g2_mux2_1 _12359_ (.A0(net617),
    .A1(net618),
    .S(net582),
    .X(_06350_));
 sg13g2_nand2_1 _12360_ (.Y(_06351_),
    .A(net593),
    .B(_06350_));
 sg13g2_o21ai_1 _12361_ (.B1(_06351_),
    .Y(_06352_),
    .A1(net593),
    .A2(_06328_));
 sg13g2_nor2_1 _12362_ (.A(net371),
    .B(_06249_),
    .Y(_06353_));
 sg13g2_a22oi_1 _12363_ (.Y(_06354_),
    .B1(_06353_),
    .B2(net393),
    .A2(_06352_),
    .A1(net369));
 sg13g2_nor2_1 _12364_ (.A(_06349_),
    .B(_06354_),
    .Y(_06355_));
 sg13g2_a22oi_1 _12365_ (.Y(_06356_),
    .B1(_04391_),
    .B2(net627),
    .A2(net341),
    .A1(net580));
 sg13g2_a22oi_1 _12366_ (.Y(_06357_),
    .B1(_06356_),
    .B2(net347),
    .A2(_06121_),
    .A1(net341));
 sg13g2_nor2_1 _12367_ (.A(net823),
    .B(_06357_),
    .Y(_06358_));
 sg13g2_a21oi_1 _12368_ (.A1(net347),
    .A2(_06355_),
    .Y(_06359_),
    .B1(_06358_));
 sg13g2_nor2_1 _12369_ (.A(net374),
    .B(_05944_),
    .Y(_06360_));
 sg13g2_a22oi_1 _12370_ (.Y(_06361_),
    .B1(_06360_),
    .B2(net363),
    .A2(_05951_),
    .A1(net372));
 sg13g2_a22oi_1 _12371_ (.Y(_06362_),
    .B1(_06361_),
    .B2(_05912_),
    .A2(_06110_),
    .A1(net367));
 sg13g2_nor3_1 _12372_ (.A(net838),
    .B(_06359_),
    .C(_06362_),
    .Y(_06363_));
 sg13g2_nand2_1 _12373_ (.Y(_06364_),
    .A(_05180_),
    .B(net618));
 sg13g2_inv_1 _12374_ (.Y(_06365_),
    .A(_06364_));
 sg13g2_nor2_1 _12375_ (.A(net847),
    .B(_05182_),
    .Y(_06366_));
 sg13g2_a21oi_1 _12376_ (.A1(net852),
    .A2(_06365_),
    .Y(_06367_),
    .B1(_06366_));
 sg13g2_nor2_1 _12377_ (.A(net564),
    .B(_06367_),
    .Y(_06368_));
 sg13g2_a21oi_1 _12378_ (.A1(net822),
    .A2(_04885_),
    .Y(_06369_),
    .B1(_06368_));
 sg13g2_nand2b_1 _12379_ (.Y(_06370_),
    .B(_06369_),
    .A_N(_06363_));
 sg13g2_a21o_1 _12380_ (.A2(_06348_),
    .A1(net339),
    .B1(_06370_),
    .X(net71));
 sg13g2_nand2_1 _12381_ (.Y(_06371_),
    .A(_06020_),
    .B(_05194_));
 sg13g2_o21ai_1 _12382_ (.B1(_06371_),
    .Y(_06372_),
    .A1(net822),
    .A2(_05179_));
 sg13g2_mux2_1 _12383_ (.A0(_05177_),
    .A1(_04928_),
    .S(net576),
    .X(_06373_));
 sg13g2_mux2_1 _12384_ (.A0(_06350_),
    .A1(_06373_),
    .S(net595),
    .X(_06374_));
 sg13g2_nand2_1 _12385_ (.Y(_06375_),
    .A(net372),
    .B(_06374_));
 sg13g2_o21ai_1 _12386_ (.B1(_06375_),
    .Y(_06376_),
    .A1(net372),
    .A2(_06262_));
 sg13g2_nor2_1 _12387_ (.A(net396),
    .B(_06376_),
    .Y(_06377_));
 sg13g2_a21oi_1 _12388_ (.A1(net396),
    .A2(_06159_),
    .Y(_06378_),
    .B1(_06377_));
 sg13g2_nor2_1 _12389_ (.A(net342),
    .B(_05999_),
    .Y(_06379_));
 sg13g2_o21ai_1 _12390_ (.B1(_06007_),
    .Y(_06380_),
    .A1(net349),
    .A2(_06379_));
 sg13g2_nor2_1 _12391_ (.A(net364),
    .B(_06163_),
    .Y(_06381_));
 sg13g2_nor2_1 _12392_ (.A(net374),
    .B(_05994_),
    .Y(_06382_));
 sg13g2_a22oi_1 _12393_ (.Y(_06383_),
    .B1(_06382_),
    .B2(net397),
    .A2(_05980_),
    .A1(net374));
 sg13g2_nor3_1 _12394_ (.A(net607),
    .B(_06381_),
    .C(_06383_),
    .Y(_06384_));
 sg13g2_a21oi_1 _12395_ (.A1(net343),
    .A2(_06380_),
    .Y(_06385_),
    .B1(_06384_));
 sg13g2_a21o_1 _12396_ (.A2(_06378_),
    .A1(net358),
    .B1(_06385_),
    .X(_06386_));
 sg13g2_a21oi_1 _12397_ (.A1(_05182_),
    .A2(net339),
    .Y(_06387_),
    .B1(net822));
 sg13g2_a21oi_1 _12398_ (.A1(_06365_),
    .A2(net339),
    .Y(_06388_),
    .B1(_04838_));
 sg13g2_a21oi_1 _12399_ (.A1(_04838_),
    .A2(_06387_),
    .Y(_06389_),
    .B1(_06388_));
 sg13g2_a221oi_1 _12400_ (.B2(net834),
    .C1(_06389_),
    .B1(_06386_),
    .A1(net638),
    .Y(_06390_),
    .A2(_06372_));
 sg13g2_or3_1 _12401_ (.A(_05182_),
    .B(_04838_),
    .C(net340),
    .X(_06391_));
 sg13g2_nand3_1 _12402_ (.B(_06364_),
    .C(net339),
    .A(_04838_),
    .Y(_06392_));
 sg13g2_mux2_1 _12403_ (.A0(_06391_),
    .A1(_06392_),
    .S(_06347_),
    .X(_06393_));
 sg13g2_nand2_1 _12404_ (.Y(net72),
    .A(_06390_),
    .B(_06393_));
 sg13g2_buf_2 fanout477 (.A(_08470_),
    .X(net477));
 sg13g2_o21ai_1 _12406_ (.B1(_06289_),
    .Y(_06395_),
    .A1(net607),
    .A2(_05888_));
 sg13g2_o21ai_1 _12407_ (.B1(_06395_),
    .Y(_06396_),
    .A1(net606),
    .A2(_05741_));
 sg13g2_mux2_1 _12408_ (.A0(_05835_),
    .A1(net618),
    .S(net576),
    .X(_06397_));
 sg13g2_mux2_1 _12409_ (.A0(_06373_),
    .A1(_06397_),
    .S(net595),
    .X(_06398_));
 sg13g2_mux2_1 _12410_ (.A0(_06283_),
    .A1(_06398_),
    .S(net373),
    .X(_06399_));
 sg13g2_mux2_1 _12411_ (.A0(_06195_),
    .A1(_06399_),
    .S(net362),
    .X(_06400_));
 sg13g2_nor4_1 _12412_ (.A(net352),
    .B(net868),
    .C(_05791_),
    .D(net342),
    .Y(_06401_));
 sg13g2_a22oi_1 _12413_ (.Y(_06402_),
    .B1(_06401_),
    .B2(net836),
    .A2(_06400_),
    .A1(net358));
 sg13g2_and2_1 _12414_ (.A(_06396_),
    .B(_06402_),
    .X(_06403_));
 sg13g2_and4_1 _12415_ (.A(_04980_),
    .B(_05242_),
    .C(_05423_),
    .D(_05430_),
    .X(_06404_));
 sg13g2_o21ai_1 _12416_ (.B1(_06404_),
    .Y(_06405_),
    .A1(_05566_),
    .A2(_05665_));
 sg13g2_a221oi_1 _12417_ (.B2(_05433_),
    .C1(_05196_),
    .B1(_05243_),
    .A1(_04980_),
    .Y(_06406_),
    .A2(_05175_));
 sg13g2_nand2_1 _12418_ (.Y(_06407_),
    .A(_06405_),
    .B(_06406_));
 sg13g2_xnor2_1 _12419_ (.Y(_06408_),
    .A(_04554_),
    .B(_06407_));
 sg13g2_a21oi_1 _12420_ (.A1(net849),
    .A2(_05835_),
    .Y(_06409_),
    .B1(net815));
 sg13g2_nand2_1 _12421_ (.Y(_06410_),
    .A(net815),
    .B(_05835_));
 sg13g2_o21ai_1 _12422_ (.B1(_06410_),
    .Y(_06411_),
    .A1(_04507_),
    .A2(_06409_));
 sg13g2_a221oi_1 _12423_ (.B2(net638),
    .C1(net831),
    .B1(_06411_),
    .A1(net819),
    .Y(_06412_),
    .A2(_04554_));
 sg13g2_o21ai_1 _12424_ (.B1(_06412_),
    .Y(_06413_),
    .A1(net356),
    .A2(_06408_));
 sg13g2_nor2b_1 _12425_ (.A(_06403_),
    .B_N(_06413_),
    .Y(net73));
 sg13g2_inv_1 _12426_ (.Y(_06414_),
    .A(net343));
 sg13g2_nand3_1 _12427_ (.B(_05863_),
    .C(_05874_),
    .A(net350),
    .Y(_06415_));
 sg13g2_a21o_1 _12428_ (.A2(_05890_),
    .A1(net350),
    .B1(net838),
    .X(_06416_));
 sg13g2_and2_1 _12429_ (.A(net367),
    .B(_06330_),
    .X(_06417_));
 sg13g2_a22oi_1 _12430_ (.Y(_06418_),
    .B1(_06417_),
    .B2(net372),
    .A2(_06087_),
    .A1(net396));
 sg13g2_mux2_1 _12431_ (.A0(_04427_),
    .A1(_05177_),
    .S(net576),
    .X(_06419_));
 sg13g2_mux2_1 _12432_ (.A0(_06397_),
    .A1(_06419_),
    .S(net595),
    .X(_06420_));
 sg13g2_nor2_1 _12433_ (.A(net362),
    .B(_06203_),
    .Y(_06421_));
 sg13g2_a22oi_1 _12434_ (.Y(_06422_),
    .B1(_06421_),
    .B2(net384),
    .A2(_06420_),
    .A1(net362));
 sg13g2_nor3_1 _12435_ (.A(net608),
    .B(_06418_),
    .C(_06422_),
    .Y(_06423_));
 sg13g2_a21oi_1 _12436_ (.A1(net609),
    .A2(_05823_),
    .Y(_06424_),
    .B1(_06423_));
 sg13g2_nor2_1 _12437_ (.A(net869),
    .B(_06424_),
    .Y(_06425_));
 sg13g2_a22oi_1 _12438_ (.Y(_06426_),
    .B1(_06416_),
    .B2(_06425_),
    .A2(_06415_),
    .A1(_06414_));
 sg13g2_inv_1 _12439_ (.Y(_06427_),
    .A(_04553_));
 sg13g2_o21ai_1 _12440_ (.B1(_06427_),
    .Y(_06428_),
    .A1(_04552_),
    .A2(_06407_));
 sg13g2_buf_2 fanout476 (.A(net477),
    .X(net476));
 sg13g2_xnor2_1 _12442_ (.Y(_06430_),
    .A(_04443_),
    .B(_06428_));
 sg13g2_a21oi_1 _12443_ (.A1(net849),
    .A2(_04427_),
    .Y(_06431_),
    .B1(net815));
 sg13g2_nand2_1 _12444_ (.Y(_06432_),
    .A(net815),
    .B(_04427_));
 sg13g2_o21ai_1 _12445_ (.B1(_06432_),
    .Y(_06433_),
    .A1(_04442_),
    .A2(_06431_));
 sg13g2_a21o_1 _12446_ (.A2(_06433_),
    .A1(net635),
    .B1(net832),
    .X(_06434_));
 sg13g2_a221oi_1 _12447_ (.B2(_06430_),
    .C1(_06434_),
    .B1(net345),
    .A1(net819),
    .Y(_06435_),
    .A2(_04443_));
 sg13g2_nor2_1 _12448_ (.A(_06426_),
    .B(_06435_),
    .Y(net74));
 sg13g2_o21ai_1 _12449_ (.B1(net625),
    .Y(_06436_),
    .A1(_04493_),
    .A2(_04496_));
 sg13g2_buf_2 fanout475 (.A(_08474_),
    .X(net475));
 sg13g2_nand2_1 _12451_ (.Y(_06438_),
    .A(_05206_),
    .B(_06436_));
 sg13g2_nand2_1 _12452_ (.Y(_06439_),
    .A(_06438_),
    .B(_05200_));
 sg13g2_or2_1 _12453_ (.X(_06440_),
    .B(_05201_),
    .A(_06438_));
 sg13g2_mux2_1 _12454_ (.A0(_06439_),
    .A1(_06440_),
    .S(_06428_),
    .X(_06441_));
 sg13g2_nand2_1 _12455_ (.Y(_06442_),
    .A(_06438_),
    .B(_05201_));
 sg13g2_o21ai_1 _12456_ (.B1(_06442_),
    .Y(_06443_),
    .A1(_06438_),
    .A2(_05200_));
 sg13g2_nor2_1 _12457_ (.A(net844),
    .B(_04503_),
    .Y(_06444_));
 sg13g2_a21oi_1 _12458_ (.A1(net849),
    .A2(_04497_),
    .Y(_06445_),
    .B1(_06444_));
 sg13g2_nand2_1 _12459_ (.Y(_06446_),
    .A(net819),
    .B(_04504_));
 sg13g2_o21ai_1 _12460_ (.B1(_06446_),
    .Y(_06447_),
    .A1(net565),
    .A2(_06445_));
 sg13g2_a21oi_1 _12461_ (.A1(net345),
    .A2(_06443_),
    .Y(_06448_),
    .B1(_06447_));
 sg13g2_o21ai_1 _12462_ (.B1(_06448_),
    .Y(_06449_),
    .A1(net356),
    .A2(_06441_));
 sg13g2_o21ai_1 _12463_ (.B1(net343),
    .Y(_06450_),
    .A1(net868),
    .A2(_05938_));
 sg13g2_o21ai_1 _12464_ (.B1(_06450_),
    .Y(_06451_),
    .A1(net608),
    .A2(_05963_));
 sg13g2_mux4_1 _12465_ (.S0(_05599_),
    .A0(_05198_),
    .A1(net624),
    .A2(_04830_),
    .A3(_04550_),
    .S1(net571),
    .X(_06452_));
 sg13g2_mux2_1 _12466_ (.A0(_06249_),
    .A1(_06452_),
    .S(net360),
    .X(_06453_));
 sg13g2_and2_1 _12467_ (.A(net396),
    .B(_06112_),
    .X(_06454_));
 sg13g2_a22oi_1 _12468_ (.Y(_06455_),
    .B1(_06454_),
    .B2(net372),
    .A2(_06352_),
    .A1(net363));
 sg13g2_a22oi_1 _12469_ (.Y(_06456_),
    .B1(_06455_),
    .B2(net868),
    .A2(_06453_),
    .A1(net374));
 sg13g2_o21ai_1 _12470_ (.B1(net352),
    .Y(_06457_),
    .A1(_05955_),
    .A2(_06456_));
 sg13g2_a21oi_1 _12471_ (.A1(_06451_),
    .A2(_06457_),
    .Y(_06458_),
    .B1(net838));
 sg13g2_a21o_1 _12472_ (.A2(_06449_),
    .A1(net840),
    .B1(_06458_),
    .X(net75));
 sg13g2_or3_1 _12473_ (.A(net607),
    .B(_05998_),
    .C(_06010_),
    .X(_06459_));
 sg13g2_mux4_1 _12474_ (.S0(net642),
    .A0(_04427_),
    .A1(_05835_),
    .A2(net612),
    .A3(_04502_),
    .S1(net581),
    .X(_06460_));
 sg13g2_mux2_1 _12475_ (.A0(_06374_),
    .A1(_06460_),
    .S(net373),
    .X(_06461_));
 sg13g2_nor2_1 _12476_ (.A(net363),
    .B(_06263_),
    .Y(_06462_));
 sg13g2_a22oi_1 _12477_ (.Y(_06463_),
    .B1(_06462_),
    .B2(net608),
    .A2(_06461_),
    .A1(net363));
 sg13g2_a22oi_1 _12478_ (.Y(_06464_),
    .B1(_06463_),
    .B2(net868),
    .A2(_06017_),
    .A1(net606));
 sg13g2_o21ai_1 _12479_ (.B1(net831),
    .Y(_06465_),
    .A1(net607),
    .A2(_06008_));
 sg13g2_a22oi_1 _12480_ (.Y(_06466_),
    .B1(_06464_),
    .B2(_06465_),
    .A2(_06459_),
    .A1(_06414_));
 sg13g2_nand2b_1 _12481_ (.Y(_06467_),
    .B(_05200_),
    .A_N(_06428_));
 sg13g2_inv_1 _12482_ (.Y(_06468_),
    .A(_04598_));
 sg13g2_nor4_1 _12483_ (.A(_04497_),
    .B(_06468_),
    .C(_05201_),
    .D(net356),
    .Y(_06469_));
 sg13g2_a22oi_1 _12484_ (.Y(_06470_),
    .B1(_04598_),
    .B2(_04497_),
    .A2(_05201_),
    .A1(_06436_));
 sg13g2_a22oi_1 _12485_ (.Y(_06471_),
    .B1(net356),
    .B2(_06470_),
    .A2(_04598_),
    .A1(_06436_));
 sg13g2_o21ai_1 _12486_ (.B1(net844),
    .Y(_06472_),
    .A1(net819),
    .A2(net623));
 sg13g2_nand2_1 _12487_ (.Y(_06473_),
    .A(_04597_),
    .B(_06472_));
 sg13g2_o21ai_1 _12488_ (.B1(_06473_),
    .Y(_06474_),
    .A1(net844),
    .A2(net623));
 sg13g2_a221oi_1 _12489_ (.B2(net635),
    .C1(net831),
    .B1(_06474_),
    .A1(net819),
    .Y(_06475_),
    .A2(_04598_));
 sg13g2_nand2b_1 _12490_ (.Y(_06476_),
    .B(_06475_),
    .A_N(_06471_));
 sg13g2_nand3_1 _12491_ (.B(_05200_),
    .C(net345),
    .A(_06436_),
    .Y(_06477_));
 sg13g2_nor3_1 _12492_ (.A(_04598_),
    .B(_06428_),
    .C(_06477_),
    .Y(_06478_));
 sg13g2_a22oi_1 _12493_ (.Y(_06479_),
    .B1(_06476_),
    .B2(_06478_),
    .A2(_06469_),
    .A1(_06467_));
 sg13g2_nor2_1 _12494_ (.A(_06466_),
    .B(_06479_),
    .Y(net76));
 sg13g2_o21ai_1 _12495_ (.B1(_06064_),
    .Y(_06480_),
    .A1(net606),
    .A2(_06066_));
 sg13g2_nor2_1 _12496_ (.A(_06096_),
    .B(_05738_),
    .Y(_06481_));
 sg13g2_o21ai_1 _12497_ (.B1(_06395_),
    .Y(_06482_),
    .A1(_06069_),
    .A2(_06481_));
 sg13g2_o21ai_1 _12498_ (.B1(_05922_),
    .Y(_06483_),
    .A1(net612),
    .A2(net571));
 sg13g2_mux2_1 _12499_ (.A0(net624),
    .A1(net620),
    .S(net581),
    .X(_06484_));
 sg13g2_mux2_1 _12500_ (.A0(_06483_),
    .A1(_06484_),
    .S(net590),
    .X(_06485_));
 sg13g2_nand2_1 _12501_ (.Y(_06486_),
    .A(net383),
    .B(_06398_));
 sg13g2_o21ai_1 _12502_ (.B1(_06486_),
    .Y(_06487_),
    .A1(net383),
    .A2(_06485_));
 sg13g2_nor2_1 _12503_ (.A(net395),
    .B(_06487_),
    .Y(_06488_));
 sg13g2_a22oi_1 _12504_ (.Y(_06489_),
    .B1(_06488_),
    .B2(net606),
    .A2(_06285_),
    .A1(net395));
 sg13g2_and3_1 _12505_ (.X(_06490_),
    .A(net606),
    .B(net362),
    .C(_06053_));
 sg13g2_o21ai_1 _12506_ (.B1(net826),
    .Y(_06491_),
    .A1(_06489_),
    .A2(_06490_));
 sg13g2_nand4_1 _12507_ (.B(_06480_),
    .C(_06482_),
    .A(net831),
    .Y(_06492_),
    .D(_06491_));
 sg13g2_inv_1 _12508_ (.Y(_06493_),
    .A(_04600_));
 sg13g2_o21ai_1 _12509_ (.B1(_05209_),
    .Y(_06494_),
    .A1(_04503_),
    .A2(_05202_));
 sg13g2_nor3_1 _12510_ (.A(_04503_),
    .B(_05209_),
    .C(_05202_),
    .Y(_06495_));
 sg13g2_a21o_1 _12511_ (.A2(_06494_),
    .A1(net612),
    .B1(_06495_),
    .X(_06496_));
 sg13g2_a21oi_1 _12512_ (.A1(_06493_),
    .A2(_06407_),
    .Y(_06497_),
    .B1(_06496_));
 sg13g2_xor2_1 _12513_ (.B(_06497_),
    .A(_04788_),
    .X(_06498_));
 sg13g2_o21ai_1 _12514_ (.B1(net842),
    .Y(_06499_),
    .A1(net817),
    .A2(net620));
 sg13g2_nor2_1 _12515_ (.A(net842),
    .B(net620),
    .Y(_06500_));
 sg13g2_a21oi_1 _12516_ (.A1(_04786_),
    .A2(_06499_),
    .Y(_06501_),
    .B1(_06500_));
 sg13g2_nor2_1 _12517_ (.A(net565),
    .B(_06501_),
    .Y(_06502_));
 sg13g2_a22oi_1 _12518_ (.Y(_06503_),
    .B1(net832),
    .B2(_06502_),
    .A2(_04788_),
    .A1(net817));
 sg13g2_o21ai_1 _12519_ (.B1(_06503_),
    .Y(_06504_),
    .A1(net356),
    .A2(_06498_));
 sg13g2_and2_1 _12520_ (.A(_06492_),
    .B(_06504_),
    .X(net78));
 sg13g2_nand2_1 _12521_ (.Y(_06505_),
    .A(_04736_),
    .B(_04738_));
 sg13g2_nand2_1 _12522_ (.Y(_06506_),
    .A(_06505_),
    .B(net344));
 sg13g2_nand3_1 _12523_ (.B(_04738_),
    .C(net344),
    .A(_04736_),
    .Y(_06507_));
 sg13g2_nand2_1 _12524_ (.Y(_06508_),
    .A(net620),
    .B(_05212_));
 sg13g2_nor2_1 _12525_ (.A(_04780_),
    .B(_05212_),
    .Y(_06509_));
 sg13g2_a21o_1 _12526_ (.A2(_06496_),
    .A1(_06508_),
    .B1(_06509_),
    .X(_06510_));
 sg13g2_nand2b_1 _12527_ (.Y(_06511_),
    .B(_06508_),
    .A_N(_04600_));
 sg13g2_a21o_1 _12528_ (.A2(_06406_),
    .A1(_06405_),
    .B1(_06511_),
    .X(_06512_));
 sg13g2_nor2b_1 _12529_ (.A(_06510_),
    .B_N(_06512_),
    .Y(_06513_));
 sg13g2_mux2_1 _12530_ (.A0(_06506_),
    .A1(_06507_),
    .S(_06513_),
    .X(_06514_));
 sg13g2_a21oi_1 _12531_ (.A1(net848),
    .A2(_05223_),
    .Y(_06515_),
    .B1(net815));
 sg13g2_nand2_1 _12532_ (.Y(_06516_),
    .A(net815),
    .B(_05223_));
 sg13g2_o21ai_1 _12533_ (.B1(_06516_),
    .Y(_06517_),
    .A1(_04734_),
    .A2(_06515_));
 sg13g2_nor2_1 _12534_ (.A(net848),
    .B(_06505_),
    .Y(_06518_));
 sg13g2_a22oi_1 _12535_ (.Y(_06519_),
    .B1(_06518_),
    .B2(net832),
    .A2(_06517_),
    .A1(net635));
 sg13g2_nand2_1 _12536_ (.Y(_06520_),
    .A(net612),
    .B(net569));
 sg13g2_o21ai_1 _12537_ (.B1(_06520_),
    .Y(_06521_),
    .A1(_04725_),
    .A2(net569));
 sg13g2_nand2_1 _12538_ (.Y(_06522_),
    .A(net640),
    .B(_06484_));
 sg13g2_o21ai_1 _12539_ (.B1(_06522_),
    .Y(_06523_),
    .A1(net640),
    .A2(_06521_));
 sg13g2_nand2_1 _12540_ (.Y(_06524_),
    .A(net369),
    .B(_06523_));
 sg13g2_o21ai_1 _12541_ (.B1(_06524_),
    .Y(_06525_),
    .A1(net369),
    .A2(_06420_));
 sg13g2_mux2_1 _12542_ (.A0(_06332_),
    .A1(_06525_),
    .S(net359),
    .X(_06526_));
 sg13g2_nand3_1 _12543_ (.B(net360),
    .C(_06088_),
    .A(net605),
    .Y(_06527_));
 sg13g2_o21ai_1 _12544_ (.B1(_06527_),
    .Y(_06528_),
    .A1(net605),
    .A2(_06526_));
 sg13g2_nor2_2 _12545_ (.A(net610),
    .B(_05888_),
    .Y(_06529_));
 sg13g2_a21o_1 _12546_ (.A2(_06529_),
    .A1(_06100_),
    .B1(net835),
    .X(_06530_));
 sg13g2_a21oi_1 _12547_ (.A1(net353),
    .A2(_06103_),
    .Y(_06531_),
    .B1(net343));
 sg13g2_a22oi_1 _12548_ (.Y(_06532_),
    .B1(_06530_),
    .B2(_06531_),
    .A2(_06528_),
    .A1(net823));
 sg13g2_a21oi_1 _12549_ (.A1(_06514_),
    .A2(_06519_),
    .Y(net79),
    .B1(_06532_));
 sg13g2_and3_1 _12550_ (.X(_06533_),
    .A(net605),
    .B(net359),
    .C(_06113_));
 sg13g2_mux2_1 _12551_ (.A0(net621),
    .A1(_05225_),
    .S(net569),
    .X(_06534_));
 sg13g2_mux2_1 _12552_ (.A0(_06521_),
    .A1(_06534_),
    .S(net589),
    .X(_06535_));
 sg13g2_mux2_1 _12553_ (.A0(_06352_),
    .A1(_06535_),
    .S(net359),
    .X(_06536_));
 sg13g2_nor2_1 _12554_ (.A(net379),
    .B(_06536_),
    .Y(_06537_));
 sg13g2_a22oi_1 _12555_ (.Y(_06538_),
    .B1(_06537_),
    .B2(net605),
    .A2(_06453_),
    .A1(net380));
 sg13g2_o21ai_1 _12556_ (.B1(net823),
    .Y(_06539_),
    .A1(_06533_),
    .A2(_06538_));
 sg13g2_a22oi_1 _12557_ (.Y(_06540_),
    .B1(net607),
    .B2(_06125_),
    .A2(_06120_),
    .A1(_06119_));
 sg13g2_nor2_1 _12558_ (.A(net343),
    .B(_06540_),
    .Y(_06541_));
 sg13g2_a22oi_1 _12559_ (.Y(_06542_),
    .B1(_06541_),
    .B2(net835),
    .A2(_06127_),
    .A1(net353));
 sg13g2_nand2_1 _12560_ (.Y(_06543_),
    .A(net622),
    .B(_04640_));
 sg13g2_o21ai_1 _12561_ (.B1(net815),
    .Y(_06544_),
    .A1(net622),
    .A2(_04640_));
 sg13g2_o21ai_1 _12562_ (.B1(_06544_),
    .Y(_06545_),
    .A1(net818),
    .A2(_06543_));
 sg13g2_nor2_1 _12563_ (.A(net848),
    .B(_04642_),
    .Y(_06546_));
 sg13g2_a21oi_1 _12564_ (.A1(net634),
    .A2(_06545_),
    .Y(_06547_),
    .B1(_06546_));
 sg13g2_nand2_1 _12565_ (.Y(_06548_),
    .A(_04642_),
    .B(net835));
 sg13g2_o21ai_1 _12566_ (.B1(net344),
    .Y(_06549_),
    .A1(_04736_),
    .A2(_06548_));
 sg13g2_and2_1 _12567_ (.A(_06547_),
    .B(_06549_),
    .X(_06550_));
 sg13g2_a21oi_1 _12568_ (.A1(_06539_),
    .A2(_06542_),
    .Y(_06551_),
    .B1(_06550_));
 sg13g2_nand3_1 _12569_ (.B(net835),
    .C(_06547_),
    .A(_04642_),
    .Y(_06552_));
 sg13g2_xnor2_1 _12570_ (.Y(_06553_),
    .A(_05949_),
    .B(_04640_));
 sg13g2_and2_1 _12571_ (.A(_06553_),
    .B(_04736_),
    .X(_06554_));
 sg13g2_nand3_1 _12572_ (.B(_06547_),
    .C(_06554_),
    .A(net835),
    .Y(_06555_));
 sg13g2_nand3b_1 _12573_ (.B(_06512_),
    .C(_04738_),
    .Y(_06556_),
    .A_N(_06510_));
 sg13g2_buf_1 fanout474 (.A(net475),
    .X(net474));
 sg13g2_mux2_1 _12575_ (.A0(_06552_),
    .A1(_06555_),
    .S(_06556_),
    .X(_06558_));
 sg13g2_nand2_1 _12576_ (.Y(_06559_),
    .A(_06551_),
    .B(_06558_));
 sg13g2_inv_1 _12577_ (.Y(net80),
    .A(_06559_));
 sg13g2_inv_1 _12578_ (.Y(_06560_),
    .A(_04689_));
 sg13g2_nor3_1 _12579_ (.A(net818),
    .B(_05215_),
    .C(_06560_),
    .Y(_06561_));
 sg13g2_a21oi_1 _12580_ (.A1(_05215_),
    .A2(_06560_),
    .Y(_06562_),
    .B1(net843));
 sg13g2_o21ai_1 _12581_ (.B1(net634),
    .Y(_06563_),
    .A1(_06561_),
    .A2(_06562_));
 sg13g2_o21ai_1 _12582_ (.B1(_06563_),
    .Y(_06564_),
    .A1(net848),
    .A2(_04690_));
 sg13g2_nor2_1 _12583_ (.A(net830),
    .B(_06564_),
    .Y(_06565_));
 sg13g2_nand3_1 _12584_ (.B(_04690_),
    .C(_06565_),
    .A(_06543_),
    .Y(_06566_));
 sg13g2_a21oi_1 _12585_ (.A1(_06556_),
    .A2(_06554_),
    .Y(_06567_),
    .B1(_06566_));
 sg13g2_and4_1 _12586_ (.A(_05222_),
    .B(_04736_),
    .C(_06556_),
    .D(_06565_),
    .X(_06568_));
 sg13g2_nor3_1 _12587_ (.A(_06543_),
    .B(_04690_),
    .C(net830),
    .Y(_06569_));
 sg13g2_nor2_1 _12588_ (.A(net355),
    .B(_06569_),
    .Y(_06570_));
 sg13g2_nor2_1 _12589_ (.A(net607),
    .B(net394),
    .Y(_06571_));
 sg13g2_nor2b_1 _12590_ (.A(_06571_),
    .B_N(net629),
    .Y(_06572_));
 sg13g2_a22oi_1 _12591_ (.Y(_06573_),
    .B1(_06572_),
    .B2(_05956_),
    .A2(_06163_),
    .A1(_06571_));
 sg13g2_nor2_1 _12592_ (.A(net394),
    .B(_06163_),
    .Y(_06574_));
 sg13g2_nor3_1 _12593_ (.A(net382),
    .B(net365),
    .C(_05999_),
    .Y(_06575_));
 sg13g2_o21ai_1 _12594_ (.B1(_06529_),
    .Y(_06576_),
    .A1(_06574_),
    .A2(_06575_));
 sg13g2_nor2b_1 _12595_ (.A(_06573_),
    .B_N(_06576_),
    .Y(_06577_));
 sg13g2_nand3_1 _12596_ (.B(net358),
    .C(_06376_),
    .A(net397),
    .Y(_06578_));
 sg13g2_mux2_1 _12597_ (.A0(_04685_),
    .A1(_05223_),
    .S(net569),
    .X(_06579_));
 sg13g2_mux2_1 _12598_ (.A0(_06534_),
    .A1(_06579_),
    .S(net588),
    .X(_06580_));
 sg13g2_mux2_1 _12599_ (.A0(_06460_),
    .A1(_06580_),
    .S(net371),
    .X(_06581_));
 sg13g2_nand2_1 _12600_ (.Y(_06582_),
    .A(net348),
    .B(_06581_));
 sg13g2_o21ai_1 _12601_ (.B1(_06582_),
    .Y(_06583_),
    .A1(net348),
    .A2(_06159_));
 sg13g2_nand3_1 _12602_ (.B(net823),
    .C(_06583_),
    .A(net360),
    .Y(_06584_));
 sg13g2_nand4_1 _12603_ (.B(_06577_),
    .C(_06578_),
    .A(net831),
    .Y(_06585_),
    .D(_06584_));
 sg13g2_o21ai_1 _12604_ (.B1(_06585_),
    .Y(_06586_),
    .A1(_06564_),
    .A2(_06570_));
 sg13g2_nor3_1 _12605_ (.A(_06567_),
    .B(_06568_),
    .C(_06586_),
    .Y(net81));
 sg13g2_mux2_1 _12606_ (.A0(_06064_),
    .A1(_06189_),
    .S(_06571_),
    .X(_06587_));
 sg13g2_nor2_1 _12607_ (.A(net621),
    .B(net581),
    .Y(_06588_));
 sg13g2_a21oi_1 _12608_ (.A1(net568),
    .A2(net578),
    .Y(_06589_),
    .B1(_06588_));
 sg13g2_nand2_1 _12609_ (.Y(_06590_),
    .A(net589),
    .B(_06589_));
 sg13g2_nand2_1 _12610_ (.Y(_06591_),
    .A(net639),
    .B(_06579_));
 sg13g2_and2_1 _12611_ (.A(_06590_),
    .B(_06591_),
    .X(_06592_));
 sg13g2_and2_1 _12612_ (.A(net380),
    .B(_06485_),
    .X(_06593_));
 sg13g2_a22oi_1 _12613_ (.Y(_06594_),
    .B1(_06593_),
    .B2(net393),
    .A2(_06592_),
    .A1(net371));
 sg13g2_a22oi_1 _12614_ (.Y(_06595_),
    .B1(_06594_),
    .B2(net606),
    .A2(_06399_),
    .A1(net395));
 sg13g2_a22oi_1 _12615_ (.Y(_06596_),
    .B1(_06595_),
    .B2(net870),
    .A2(_06197_),
    .A1(net606));
 sg13g2_nor3_1 _12616_ (.A(net836),
    .B(_06587_),
    .C(_06596_),
    .Y(_06597_));
 sg13g2_xor2_1 _12617_ (.B(_05675_),
    .A(net338),
    .X(_06598_));
 sg13g2_o21ai_1 _12618_ (.B1(net841),
    .Y(_06599_),
    .A1(net816),
    .A2(net568));
 sg13g2_nand2_1 _12619_ (.Y(_06600_),
    .A(_04060_),
    .B(_06599_));
 sg13g2_o21ai_1 _12620_ (.B1(_06600_),
    .Y(_06601_),
    .A1(net841),
    .A2(_05673_));
 sg13g2_a221oi_1 _12621_ (.B2(net634),
    .C1(net830),
    .B1(_06601_),
    .A1(net816),
    .Y(_06602_),
    .A2(_05675_));
 sg13g2_inv_1 _12622_ (.Y(_06603_),
    .A(_06602_));
 sg13g2_a21oi_1 _12623_ (.A1(net345),
    .A2(_06598_),
    .Y(_06604_),
    .B1(_06603_));
 sg13g2_nor2_1 _12624_ (.A(_06597_),
    .B(_06604_),
    .Y(net82));
 sg13g2_a21o_1 _12625_ (.A2(net338),
    .A1(_04060_),
    .B1(_04050_),
    .X(_06605_));
 sg13g2_buf_2 fanout473 (.A(net474),
    .X(net473));
 sg13g2_or2_1 _12627_ (.X(_06607_),
    .B(net338),
    .A(_04060_));
 sg13g2_buf_2 fanout472 (.A(net475),
    .X(net472));
 sg13g2_nand2_1 _12629_ (.Y(_06609_),
    .A(_06605_),
    .B(_06607_));
 sg13g2_xnor2_1 _12630_ (.Y(_06610_),
    .A(_05671_),
    .B(_06609_));
 sg13g2_nor2_1 _12631_ (.A(net369),
    .B(net359),
    .Y(_06611_));
 sg13g2_mux2_1 _12632_ (.A0(net632),
    .A1(_05215_),
    .S(net569),
    .X(_06612_));
 sg13g2_nor2_1 _12633_ (.A(net639),
    .B(_06612_),
    .Y(_06613_));
 sg13g2_a21oi_1 _12634_ (.A1(net639),
    .A2(_06589_),
    .Y(_06614_),
    .B1(_06613_));
 sg13g2_nor2_1 _12635_ (.A(net342),
    .B(_06614_),
    .Y(_06615_));
 sg13g2_nand2_1 _12636_ (.Y(_06616_),
    .A(net379),
    .B(net359));
 sg13g2_nand2_1 _12637_ (.Y(_06617_),
    .A(_06070_),
    .B(_06420_));
 sg13g2_o21ai_1 _12638_ (.B1(_06617_),
    .Y(_06618_),
    .A1(_06616_),
    .A2(_06523_));
 sg13g2_a22oi_1 _12639_ (.Y(_06619_),
    .B1(_06615_),
    .B2(_06618_),
    .A2(_06330_),
    .A1(_06611_));
 sg13g2_nand3_1 _12640_ (.B(_05886_),
    .C(_06529_),
    .A(net361),
    .Y(_06620_));
 sg13g2_o21ai_1 _12641_ (.B1(_06620_),
    .Y(_06621_),
    .A1(_05790_),
    .A2(_06619_));
 sg13g2_nand2b_1 _12642_ (.Y(_06622_),
    .B(_05853_),
    .A_N(_06213_));
 sg13g2_a21oi_1 _12643_ (.A1(net825),
    .A2(_06207_),
    .Y(_06623_),
    .B1(_06414_));
 sg13g2_a22oi_1 _12644_ (.Y(_06624_),
    .B1(_06623_),
    .B2(net836),
    .A2(_06622_),
    .A1(net350));
 sg13g2_inv_1 _12645_ (.Y(_06625_),
    .A(_04110_));
 sg13g2_nor3_1 _12646_ (.A(net818),
    .B(net633),
    .C(_06625_),
    .Y(_06626_));
 sg13g2_nor2_1 _12647_ (.A(net843),
    .B(_04112_),
    .Y(_06627_));
 sg13g2_o21ai_1 _12648_ (.B1(net634),
    .Y(_06628_),
    .A1(_06626_),
    .A2(_06627_));
 sg13g2_o21ai_1 _12649_ (.B1(_06628_),
    .Y(_06629_),
    .A1(net848),
    .A2(_05671_));
 sg13g2_a22oi_1 _12650_ (.Y(_06630_),
    .B1(_06624_),
    .B2(_06629_),
    .A2(_06621_),
    .A1(net830));
 sg13g2_buf_2 fanout471 (.A(net475),
    .X(net471));
 sg13g2_o21ai_1 _12652_ (.B1(_06630_),
    .Y(net83),
    .A1(net340),
    .A2(_06610_));
 sg13g2_nor3_1 _12653_ (.A(_04113_),
    .B(_05677_),
    .C(net340),
    .Y(_06632_));
 sg13g2_xnor2_1 _12654_ (.Y(_06633_),
    .A(_05942_),
    .B(_04173_));
 sg13g2_nor3_1 _12655_ (.A(_05676_),
    .B(_06633_),
    .C(net340),
    .Y(_06634_));
 sg13g2_mux2_1 _12656_ (.A0(_06632_),
    .A1(_06634_),
    .S(net338),
    .X(_06635_));
 sg13g2_nand2_1 _12657_ (.Y(_06636_),
    .A(net350),
    .B(_06245_));
 sg13g2_nor3_1 _12658_ (.A(net351),
    .B(net869),
    .C(_06252_),
    .Y(_06637_));
 sg13g2_mux2_1 _12659_ (.A0(net631),
    .A1(net568),
    .S(net569),
    .X(_06638_));
 sg13g2_mux2_1 _12660_ (.A0(_06612_),
    .A1(_06638_),
    .S(net588),
    .X(_06639_));
 sg13g2_mux2_1 _12661_ (.A0(_06452_),
    .A1(_06639_),
    .S(net359),
    .X(_06640_));
 sg13g2_nor2_1 _12662_ (.A(net379),
    .B(_06640_),
    .Y(_06641_));
 sg13g2_a21oi_1 _12663_ (.A1(net380),
    .A2(_06536_),
    .Y(_06642_),
    .B1(_06641_));
 sg13g2_nand2_1 _12664_ (.Y(_06643_),
    .A(net361),
    .B(_06529_));
 sg13g2_nand2b_1 _12665_ (.Y(_06644_),
    .B(_05947_),
    .A_N(_06643_));
 sg13g2_o21ai_1 _12666_ (.B1(_06644_),
    .Y(_06645_),
    .A1(_05790_),
    .A2(_06642_));
 sg13g2_a22oi_1 _12667_ (.Y(_06646_),
    .B1(_06637_),
    .B2(_06645_),
    .A2(_06636_),
    .A1(_06414_));
 sg13g2_nor3_1 _12668_ (.A(net816),
    .B(net631),
    .C(_04173_),
    .Y(_06647_));
 sg13g2_a21oi_1 _12669_ (.A1(net815),
    .A2(_04179_),
    .Y(_06648_),
    .B1(_06647_));
 sg13g2_nand3_1 _12670_ (.B(_05677_),
    .C(_06141_),
    .A(_04113_),
    .Y(_06649_));
 sg13g2_o21ai_1 _12671_ (.B1(_06649_),
    .Y(_06650_),
    .A1(net565),
    .A2(_06648_));
 sg13g2_nor2b_1 _12672_ (.A(_05671_),
    .B_N(_05675_),
    .Y(_06651_));
 sg13g2_nor3_1 _12673_ (.A(_04113_),
    .B(_06651_),
    .C(net340),
    .Y(_06652_));
 sg13g2_o21ai_1 _12674_ (.B1(_06633_),
    .Y(_06653_),
    .A1(net816),
    .A2(_06652_));
 sg13g2_nor2b_1 _12675_ (.A(_06650_),
    .B_N(_06653_),
    .Y(_06654_));
 sg13g2_o21ai_1 _12676_ (.B1(_06654_),
    .Y(_06655_),
    .A1(net837),
    .A2(_06646_));
 sg13g2_nor2_1 _12677_ (.A(_06635_),
    .B(_06655_),
    .Y(_06656_));
 sg13g2_inv_1 _12678_ (.Y(net84),
    .A(_06656_));
 sg13g2_and4_1 _12679_ (.A(_04179_),
    .B(_06651_),
    .C(_05678_),
    .D(net344),
    .X(_06657_));
 sg13g2_o21ai_1 _12680_ (.B1(_05678_),
    .Y(_06658_),
    .A1(_04113_),
    .A2(_04175_));
 sg13g2_mux2_1 _12681_ (.A0(_05678_),
    .A1(_06658_),
    .S(_04179_),
    .X(_06659_));
 sg13g2_o21ai_1 _12682_ (.B1(net843),
    .Y(_06660_),
    .A1(net818),
    .A2(_03989_));
 sg13g2_nand2_1 _12683_ (.Y(_06661_),
    .A(_03901_),
    .B(_06660_));
 sg13g2_o21ai_1 _12684_ (.B1(_06661_),
    .Y(_06662_),
    .A1(net841),
    .A2(_03989_));
 sg13g2_nor2_1 _12685_ (.A(net848),
    .B(_05678_),
    .Y(_06663_));
 sg13g2_a22oi_1 _12686_ (.Y(_06664_),
    .B1(_06663_),
    .B2(net830),
    .A2(_06662_),
    .A1(net635));
 sg13g2_o21ai_1 _12687_ (.B1(_06664_),
    .Y(_06665_),
    .A1(net355),
    .A2(_06659_));
 sg13g2_a21oi_1 _12688_ (.A1(net338),
    .A2(_06657_),
    .Y(_06666_),
    .B1(_06665_));
 sg13g2_nand2_1 _12689_ (.Y(_06667_),
    .A(net338),
    .B(_06651_));
 sg13g2_nor3_1 _12690_ (.A(_04113_),
    .B(_04175_),
    .C(_05678_),
    .Y(_06668_));
 sg13g2_nand3_1 _12691_ (.B(net344),
    .C(_06668_),
    .A(_06667_),
    .Y(_06669_));
 sg13g2_nand2_1 _12692_ (.Y(_06670_),
    .A(net347),
    .B(net341));
 sg13g2_nor2_1 _12693_ (.A(_06001_),
    .B(_06670_),
    .Y(_06671_));
 sg13g2_a22oi_1 _12694_ (.Y(_06672_),
    .B1(_06671_),
    .B2(_05956_),
    .A2(_06670_),
    .A1(net629));
 sg13g2_o21ai_1 _12695_ (.B1(net831),
    .Y(_06673_),
    .A1(_06004_),
    .A2(_06643_));
 sg13g2_nor2_1 _12696_ (.A(net632),
    .B(net578),
    .Y(_06674_));
 sg13g2_a21oi_1 _12697_ (.A1(_04177_),
    .A2(net578),
    .Y(_06675_),
    .B1(_06674_));
 sg13g2_mux2_1 _12698_ (.A0(_06638_),
    .A1(_06675_),
    .S(net588),
    .X(_06676_));
 sg13g2_nor2_1 _12699_ (.A(net369),
    .B(_06580_),
    .Y(_06677_));
 sg13g2_a22oi_1 _12700_ (.Y(_06678_),
    .B1(_06677_),
    .B2(net392),
    .A2(_06676_),
    .A1(net369));
 sg13g2_a22oi_1 _12701_ (.Y(_06679_),
    .B1(_06678_),
    .B2(net605),
    .A2(_06461_),
    .A1(net392));
 sg13g2_a22oi_1 _12702_ (.Y(_06680_),
    .B1(_06679_),
    .B2(net870),
    .A2(_06265_),
    .A1(net605));
 sg13g2_nor3_1 _12703_ (.A(_06672_),
    .B(_06673_),
    .C(_06680_),
    .Y(_06681_));
 sg13g2_a21oi_1 _12704_ (.A1(_06666_),
    .A2(_06669_),
    .Y(net85),
    .B1(_06681_));
 sg13g2_o21ai_1 _12705_ (.B1(net841),
    .Y(_06682_),
    .A1(_05735_),
    .A2(net816));
 sg13g2_nand2_1 _12706_ (.Y(_06683_),
    .A(_04285_),
    .B(_06682_));
 sg13g2_o21ai_1 _12707_ (.B1(_06683_),
    .Y(_06684_),
    .A1(_05735_),
    .A2(net841));
 sg13g2_a221oi_1 _12708_ (.B2(net634),
    .C1(net830),
    .B1(_06684_),
    .A1(net816),
    .Y(_06685_),
    .A2(_04288_));
 sg13g2_a21oi_1 _12709_ (.A1(net338),
    .A2(_05680_),
    .Y(_06686_),
    .B1(_04183_));
 sg13g2_xnor2_1 _12710_ (.Y(_06687_),
    .A(_04288_),
    .B(_06686_));
 sg13g2_nand2_1 _12711_ (.Y(_06688_),
    .A(net344),
    .B(_06687_));
 sg13g2_nor2_1 _12712_ (.A(net348),
    .B(_06287_),
    .Y(_06689_));
 sg13g2_nor2_1 _12713_ (.A(net588),
    .B(_06675_),
    .Y(_06690_));
 sg13g2_nand2_1 _12714_ (.Y(_06691_),
    .A(_05735_),
    .B(net578));
 sg13g2_o21ai_1 _12715_ (.B1(_06691_),
    .Y(_06692_),
    .A1(_05942_),
    .A2(net578));
 sg13g2_nor2_1 _12716_ (.A(net639),
    .B(_06692_),
    .Y(_06693_));
 sg13g2_nor3_1 _12717_ (.A(net379),
    .B(_06690_),
    .C(_06693_),
    .Y(_06694_));
 sg13g2_a22oi_1 _12718_ (.Y(_06695_),
    .B1(_06694_),
    .B2(net392),
    .A2(_06592_),
    .A1(net379));
 sg13g2_a22oi_1 _12719_ (.Y(_06696_),
    .B1(_06695_),
    .B2(net605),
    .A2(_06487_),
    .A1(net393));
 sg13g2_nor2_1 _12720_ (.A(_06689_),
    .B(_06696_),
    .Y(_06697_));
 sg13g2_mux2_1 _12721_ (.A0(_06071_),
    .A1(_06064_),
    .S(_06670_),
    .X(_06698_));
 sg13g2_a22oi_1 _12722_ (.Y(_06699_),
    .B1(_06698_),
    .B2(net836),
    .A2(_06697_),
    .A1(net823));
 sg13g2_a21oi_1 _12723_ (.A1(_06685_),
    .A2(_06688_),
    .Y(net86),
    .B1(_06699_));
 sg13g2_nor2_1 _12724_ (.A(net588),
    .B(_06692_),
    .Y(_06700_));
 sg13g2_nand2_1 _12725_ (.Y(_06701_),
    .A(_03989_),
    .B(net569));
 sg13g2_o21ai_1 _12726_ (.B1(_06701_),
    .Y(_06702_),
    .A1(_05868_),
    .A2(net569));
 sg13g2_nor2_1 _12727_ (.A(net639),
    .B(_06702_),
    .Y(_06703_));
 sg13g2_nor3_1 _12728_ (.A(net379),
    .B(_06700_),
    .C(_06703_),
    .Y(_06704_));
 sg13g2_a22oi_1 _12729_ (.Y(_06705_),
    .B1(_06704_),
    .B2(net392),
    .A2(_06614_),
    .A1(net379));
 sg13g2_nor2_1 _12730_ (.A(net359),
    .B(_06525_),
    .Y(_06706_));
 sg13g2_o21ai_1 _12731_ (.B1(net347),
    .Y(_06707_),
    .A1(_06705_),
    .A2(_06706_));
 sg13g2_o21ai_1 _12732_ (.B1(_06707_),
    .Y(_06708_),
    .A1(net347),
    .A2(_06334_));
 sg13g2_a21o_1 _12733_ (.A2(_06337_),
    .A1(net349),
    .B1(net835),
    .X(_06709_));
 sg13g2_a21oi_1 _12734_ (.A1(net349),
    .A2(_06336_),
    .Y(_06710_),
    .B1(net343));
 sg13g2_a22oi_1 _12735_ (.Y(_06711_),
    .B1(_06709_),
    .B2(_06710_),
    .A2(_06708_),
    .A1(net823));
 sg13g2_nor2b_1 _12736_ (.A(_05686_),
    .B_N(_04236_),
    .Y(_06712_));
 sg13g2_nor2b_1 _12737_ (.A(_04183_),
    .B_N(_06712_),
    .Y(_06713_));
 sg13g2_nor2_1 _12738_ (.A(_04278_),
    .B(_04285_),
    .Y(_06714_));
 sg13g2_nor2_1 _12739_ (.A(_04236_),
    .B(_06714_),
    .Y(_06715_));
 sg13g2_and2_1 _12740_ (.A(_05680_),
    .B(_06715_),
    .X(_06716_));
 sg13g2_mux2_1 _12741_ (.A0(_06713_),
    .A1(_06716_),
    .S(_05669_),
    .X(_06717_));
 sg13g2_nor2_1 _12742_ (.A(_04183_),
    .B(_05680_),
    .Y(_06718_));
 sg13g2_mux2_1 _12743_ (.A0(_05686_),
    .A1(_06714_),
    .S(_04236_),
    .X(_06719_));
 sg13g2_a221oi_1 _12744_ (.B2(_06718_),
    .C1(_06719_),
    .B1(_06712_),
    .A1(_04183_),
    .Y(_06720_),
    .A2(_06715_));
 sg13g2_nor2b_1 _12745_ (.A(_06717_),
    .B_N(_06720_),
    .Y(_06721_));
 sg13g2_o21ai_1 _12746_ (.B1(net841),
    .Y(_06722_),
    .A1(_04235_),
    .A2(net816));
 sg13g2_nand2_1 _12747_ (.Y(_06723_),
    .A(_04191_),
    .B(_06722_));
 sg13g2_o21ai_1 _12748_ (.B1(_06723_),
    .Y(_06724_),
    .A1(_04235_),
    .A2(net841));
 sg13g2_a221oi_1 _12749_ (.B2(net634),
    .C1(net832),
    .B1(_06724_),
    .A1(net816),
    .Y(_06725_),
    .A2(_04236_));
 sg13g2_o21ai_1 _12750_ (.B1(_06725_),
    .Y(_06726_),
    .A1(net355),
    .A2(_06721_));
 sg13g2_nor2b_1 _12751_ (.A(_06711_),
    .B_N(_06726_),
    .Y(net87));
 sg13g2_nor2_1 _12752_ (.A(_04278_),
    .B(net579),
    .Y(_06727_));
 sg13g2_a21oi_1 _12753_ (.A1(net626),
    .A2(net579),
    .Y(_06728_),
    .B1(_06727_));
 sg13g2_nor2_1 _12754_ (.A(net588),
    .B(_06702_),
    .Y(_06729_));
 sg13g2_a22oi_1 _12755_ (.Y(_06730_),
    .B1(_06729_),
    .B2(net342),
    .A2(_06728_),
    .A1(net588));
 sg13g2_nor2_1 _12756_ (.A(_06096_),
    .B(_06535_),
    .Y(_06731_));
 sg13g2_a22oi_1 _12757_ (.Y(_06732_),
    .B1(_06730_),
    .B2(_06731_),
    .A2(_06640_),
    .A1(net380));
 sg13g2_inv_1 _12758_ (.Y(_06733_),
    .A(_06732_));
 sg13g2_nor2_1 _12759_ (.A(net347),
    .B(_06355_),
    .Y(_06734_));
 sg13g2_a22oi_1 _12760_ (.Y(_06735_),
    .B1(_06734_),
    .B2(net870),
    .A2(_06733_),
    .A1(net347));
 sg13g2_nand2_1 _12761_ (.Y(_06736_),
    .A(net627),
    .B(net342));
 sg13g2_o21ai_1 _12762_ (.B1(_06736_),
    .Y(_06737_),
    .A1(net342),
    .A2(_05958_));
 sg13g2_a21oi_1 _12763_ (.A1(net347),
    .A2(_06737_),
    .Y(_06738_),
    .B1(net343));
 sg13g2_nor3_1 _12764_ (.A(net381),
    .B(_05940_),
    .C(_06643_),
    .Y(_06739_));
 sg13g2_nor4_2 _12765_ (.A(net835),
    .B(_06735_),
    .C(_06738_),
    .Y(_06740_),
    .D(_06739_));
 sg13g2_or2_1 _12766_ (.X(_06741_),
    .B(_05690_),
    .A(_05688_));
 sg13g2_inv_1 _12767_ (.Y(_06742_),
    .A(_05707_));
 sg13g2_nor3_1 _12768_ (.A(_06741_),
    .B(_05705_),
    .C(_06742_),
    .Y(_06743_));
 sg13g2_xor2_1 _12769_ (.B(_06743_),
    .A(_04398_),
    .X(_06744_));
 sg13g2_o21ai_1 _12770_ (.B1(net841),
    .Y(_06745_),
    .A1(net626),
    .A2(net817));
 sg13g2_nand2_1 _12771_ (.Y(_06746_),
    .A(_04396_),
    .B(_06745_));
 sg13g2_o21ai_1 _12772_ (.B1(_06746_),
    .Y(_06747_),
    .A1(net626),
    .A2(net842));
 sg13g2_a221oi_1 _12773_ (.B2(net634),
    .C1(net830),
    .B1(_06747_),
    .A1(net817),
    .Y(_06748_),
    .A2(_04398_));
 sg13g2_o21ai_1 _12774_ (.B1(_06748_),
    .Y(_06749_),
    .A1(net355),
    .A2(_06744_));
 sg13g2_nor2b_1 _12775_ (.A(_06740_),
    .B_N(_06749_),
    .Y(net89));
 sg13g2_xnor2_1 _12776_ (.Y(_06750_),
    .A(net629),
    .B(_04352_));
 sg13g2_nand3_1 _12777_ (.B(net344),
    .C(_06750_),
    .A(_05692_),
    .Y(_06751_));
 sg13g2_nor2_1 _12778_ (.A(_04289_),
    .B(_06751_),
    .Y(_06752_));
 sg13g2_nand3_1 _12779_ (.B(_05680_),
    .C(_06752_),
    .A(_05669_),
    .Y(_06753_));
 sg13g2_nand2_1 _12780_ (.Y(_06754_),
    .A(net345),
    .B(_06750_));
 sg13g2_nor2b_1 _12781_ (.A(_06754_),
    .B_N(_05694_),
    .Y(_06755_));
 sg13g2_o21ai_1 _12782_ (.B1(net842),
    .Y(_06756_),
    .A1(net817),
    .A2(net630));
 sg13g2_nand2b_1 _12783_ (.Y(_06757_),
    .B(_06756_),
    .A_N(_04352_));
 sg13g2_o21ai_1 _12784_ (.B1(_06757_),
    .Y(_06758_),
    .A1(net842),
    .A2(net629));
 sg13g2_nor3_1 _12785_ (.A(_05692_),
    .B(net356),
    .C(_06750_),
    .Y(_06759_));
 sg13g2_a22oi_1 _12786_ (.Y(_06760_),
    .B1(_06759_),
    .B2(net830),
    .A2(_06758_),
    .A1(net634));
 sg13g2_o21ai_1 _12787_ (.B1(_06760_),
    .Y(_06761_),
    .A1(net848),
    .A2(_06750_));
 sg13g2_a22oi_1 _12788_ (.Y(_06762_),
    .B1(_06755_),
    .B2(_06761_),
    .A2(_06752_),
    .A1(_04183_));
 sg13g2_and2_1 _12789_ (.A(_06753_),
    .B(_06762_),
    .X(_06763_));
 sg13g2_nor2_1 _12790_ (.A(_05705_),
    .B(_06742_),
    .Y(_06764_));
 sg13g2_a22oi_1 _12791_ (.Y(_06765_),
    .B1(net355),
    .B2(_06750_),
    .A2(_04396_),
    .A1(_05684_));
 sg13g2_nor2b_1 _12792_ (.A(_06741_),
    .B_N(_06765_),
    .Y(_06766_));
 sg13g2_nand2_1 _12793_ (.Y(_06767_),
    .A(_06764_),
    .B(_06766_));
 sg13g2_nor2_1 _12794_ (.A(net352),
    .B(_06378_),
    .Y(_06768_));
 sg13g2_nor2_1 _12795_ (.A(_05868_),
    .B(net578),
    .Y(_06769_));
 sg13g2_a22oi_1 _12796_ (.Y(_06770_),
    .B1(_06769_),
    .B2(net639),
    .A2(net578),
    .A1(net627));
 sg13g2_a22oi_1 _12797_ (.Y(_06771_),
    .B1(_06770_),
    .B2(net380),
    .A2(_06728_),
    .A1(net640));
 sg13g2_a22oi_1 _12798_ (.Y(_06772_),
    .B1(_06771_),
    .B2(net392),
    .A2(_06676_),
    .A1(net379));
 sg13g2_a22oi_1 _12799_ (.Y(_06773_),
    .B1(_06772_),
    .B2(net605),
    .A2(_06581_),
    .A1(net393));
 sg13g2_nor3_1 _12800_ (.A(net870),
    .B(_06768_),
    .C(_06773_),
    .Y(_06774_));
 sg13g2_a22oi_1 _12801_ (.Y(_06775_),
    .B1(net836),
    .B2(_06064_),
    .A2(_06529_),
    .A1(_06379_));
 sg13g2_nor2b_1 _12802_ (.A(_06774_),
    .B_N(_06775_),
    .Y(_06776_));
 sg13g2_a21oi_1 _12803_ (.A1(_06763_),
    .A2(_06767_),
    .Y(net90),
    .B1(_06776_));
 sg13g2_nor3_1 _12804_ (.A(net1250),
    .B(net1039),
    .C(net1024),
    .Y(_06777_));
 sg13g2_or2_1 _12805_ (.X(_06778_),
    .B(_06777_),
    .A(_03837_));
 sg13g2_buf_2 fanout470 (.A(net475),
    .X(net470));
 sg13g2_nor2_2 _12807_ (.A(net895),
    .B(net892),
    .Y(_06780_));
 sg13g2_buf_1 fanout469 (.A(net470),
    .X(net469));
 sg13g2_nor2_1 _12809_ (.A(_03837_),
    .B(_06777_),
    .Y(_06782_));
 sg13g2_nor2_1 _12810_ (.A(_01023_),
    .B(net885),
    .Y(_06783_));
 sg13g2_a21oi_1 _12811_ (.A1(_05641_),
    .A2(_05644_),
    .Y(_06784_),
    .B1(_05648_));
 sg13g2_a22oi_1 _12812_ (.Y(_06785_),
    .B1(_06783_),
    .B2(_06784_),
    .A2(_06780_),
    .A1(_05656_));
 sg13g2_a21o_1 _12813_ (.A2(_03839_),
    .A1(net1375),
    .B1(_03841_),
    .X(_06786_));
 sg13g2_buf_2 fanout468 (.A(net470),
    .X(net468));
 sg13g2_a21o_1 _12815_ (.A2(_05644_),
    .A1(_05641_),
    .B1(_05648_),
    .X(_06788_));
 sg13g2_nand3_1 _12816_ (.B(_03746_),
    .C(_05449_),
    .A(net939),
    .Y(_06789_));
 sg13g2_buf_1 fanout467 (.A(_02174_),
    .X(net467));
 sg13g2_nor2_1 _12818_ (.A(_06788_),
    .B(_06789_),
    .Y(_06791_));
 sg13g2_and2_1 _12819_ (.A(_06784_),
    .B(_06783_),
    .X(_06792_));
 sg13g2_a221oi_1 _12820_ (.B2(_06791_),
    .C1(_06792_),
    .B1(_05656_),
    .A1(net647),
    .Y(_06793_),
    .A2(_06786_));
 sg13g2_or2_1 _12821_ (.X(_06794_),
    .B(_06793_),
    .A(_06785_));
 sg13g2_buf_1 fanout466 (.A(net467),
    .X(net466));
 sg13g2_nand2_1 _12823_ (.Y(_06796_),
    .A(_05567_),
    .B(_05580_));
 sg13g2_nand3_1 _12824_ (.B(_05582_),
    .C(_06780_),
    .A(_05578_),
    .Y(_06797_));
 sg13g2_buf_2 fanout465 (.A(net466),
    .X(net465));
 sg13g2_nor2_1 _12826_ (.A(_01024_),
    .B(net888),
    .Y(_06799_));
 sg13g2_nand2_1 _12827_ (.Y(_06800_),
    .A(_05567_),
    .B(_06799_));
 sg13g2_o21ai_1 _12828_ (.B1(_06800_),
    .Y(_06801_),
    .A1(_06796_),
    .A2(_06797_));
 sg13g2_a22oi_1 _12829_ (.Y(_06802_),
    .B1(_06799_),
    .B2(_05567_),
    .A2(_06780_),
    .A1(_05591_));
 sg13g2_nor2_1 _12830_ (.A(_06801_),
    .B(_06802_),
    .Y(_06803_));
 sg13g2_xnor2_1 _12831_ (.Y(_06804_),
    .A(_06794_),
    .B(_06803_));
 sg13g2_inv_1 _12832_ (.Y(_06805_),
    .A(_03389_));
 sg13g2_xor2_1 _12833_ (.B(net627),
    .A(_03418_),
    .X(_06806_));
 sg13g2_o21ai_1 _12834_ (.B1(_03376_),
    .Y(_06807_),
    .A1(_04211_),
    .A2(_04233_));
 sg13g2_nor3_1 _12835_ (.A(_03359_),
    .B(_04261_),
    .C(_04276_),
    .Y(_06808_));
 sg13g2_nor3_1 _12836_ (.A(_03376_),
    .B(_04211_),
    .C(_04233_),
    .Y(_06809_));
 sg13g2_a21o_1 _12837_ (.A2(_06808_),
    .A1(_06807_),
    .B1(_06809_),
    .X(_06810_));
 sg13g2_a22oi_1 _12838_ (.Y(_06811_),
    .B1(_06806_),
    .B2(_06810_),
    .A2(net626),
    .A1(_06805_));
 sg13g2_nand2_1 _12839_ (.Y(_06812_),
    .A(_03389_),
    .B(_05684_));
 sg13g2_nor2_1 _12840_ (.A(net985),
    .B(_03814_),
    .Y(_06813_));
 sg13g2_nand4_1 _12841_ (.B(_02570_),
    .C(_03418_),
    .A(net1239),
    .Y(_06814_),
    .D(_06813_));
 sg13g2_nand3_1 _12842_ (.B(_02570_),
    .C(_06813_),
    .A(net1239),
    .Y(_06815_));
 sg13g2_nand2b_1 _12843_ (.Y(_06816_),
    .B(_06815_),
    .A_N(_03418_));
 sg13g2_mux2_1 _12844_ (.A0(_06814_),
    .A1(_06816_),
    .S(net628),
    .X(_06817_));
 sg13g2_o21ai_1 _12845_ (.B1(_06817_),
    .Y(_06818_),
    .A1(_06806_),
    .A2(_06812_));
 sg13g2_or2_1 _12846_ (.X(_06819_),
    .B(_06818_),
    .A(_06811_));
 sg13g2_buf_2 fanout464 (.A(net467),
    .X(net464));
 sg13g2_and2_1 _12848_ (.A(_03889_),
    .B(_04177_),
    .X(_06821_));
 sg13g2_a21oi_1 _12849_ (.A1(_03314_),
    .A2(_05942_),
    .Y(_06822_),
    .B1(_06821_));
 sg13g2_nand2b_1 _12850_ (.Y(_06823_),
    .B(net632),
    .A_N(_03296_));
 sg13g2_inv_1 _12851_ (.Y(_06824_),
    .A(_03264_));
 sg13g2_o21ai_1 _12852_ (.B1(_03296_),
    .Y(_06825_),
    .A1(_04079_),
    .A2(_04100_));
 sg13g2_o21ai_1 _12853_ (.B1(_06825_),
    .Y(_06826_),
    .A1(_06824_),
    .A2(net568));
 sg13g2_nand2b_1 _12854_ (.Y(_06827_),
    .B(net631),
    .A_N(_03314_));
 sg13g2_nand3_1 _12855_ (.B(_06826_),
    .C(_06827_),
    .A(_06823_),
    .Y(_06828_));
 sg13g2_nor2_1 _12856_ (.A(_03889_),
    .B(_04177_),
    .Y(_06829_));
 sg13g2_a21oi_1 _12857_ (.A1(_06822_),
    .A2(_06828_),
    .Y(_06830_),
    .B1(_06829_));
 sg13g2_o21ai_1 _12858_ (.B1(_03359_),
    .Y(_06831_),
    .A1(_04261_),
    .A2(_04276_));
 sg13g2_a21o_1 _12859_ (.A2(_06831_),
    .A1(_06807_),
    .B1(_06809_),
    .X(_06832_));
 sg13g2_a22oi_1 _12860_ (.Y(_06833_),
    .B1(_06806_),
    .B2(_06832_),
    .A2(net626),
    .A1(_06805_));
 sg13g2_or2_1 _12861_ (.X(_06834_),
    .B(_06833_),
    .A(_06818_));
 sg13g2_a21oi_1 _12862_ (.A1(_06819_),
    .A2(_06830_),
    .Y(_06835_),
    .B1(_06834_));
 sg13g2_and2_1 _12863_ (.A(_03049_),
    .B(_03177_),
    .X(_06836_));
 sg13g2_buf_2 fanout463 (.A(net467),
    .X(net463));
 sg13g2_nor2_1 _12865_ (.A(_04725_),
    .B(_06836_),
    .Y(_06838_));
 sg13g2_nor4_1 _12866_ (.A(net949),
    .B(_03155_),
    .C(_04758_),
    .D(_04778_),
    .Y(_06839_));
 sg13g2_a21oi_1 _12867_ (.A1(_04725_),
    .A2(_06836_),
    .Y(_06840_),
    .B1(_06839_));
 sg13g2_or2_1 _12868_ (.X(_06841_),
    .B(_03206_),
    .A(net949));
 sg13g2_buf_1 fanout462 (.A(net467),
    .X(net462));
 sg13g2_o21ai_1 _12870_ (.B1(_06841_),
    .Y(_06843_),
    .A1(_06838_),
    .A2(_06840_));
 sg13g2_and2_1 _12871_ (.A(_03236_),
    .B(_04685_),
    .X(_06844_));
 sg13g2_buf_2 fanout461 (.A(net462),
    .X(net461));
 sg13g2_nor2_1 _12873_ (.A(net621),
    .B(_06844_),
    .Y(_06846_));
 sg13g2_nor4_1 _12874_ (.A(_06841_),
    .B(_06844_),
    .C(_06838_),
    .D(_06840_),
    .Y(_06847_));
 sg13g2_nor2_1 _12875_ (.A(_03236_),
    .B(_04685_),
    .Y(_06848_));
 sg13g2_a22oi_1 _12876_ (.Y(_06849_),
    .B1(_06847_),
    .B2(_06848_),
    .A2(_06846_),
    .A1(_06843_));
 sg13g2_nor2_1 _12877_ (.A(net950),
    .B(_03078_),
    .Y(_06850_));
 sg13g2_o21ai_1 _12878_ (.B1(net623),
    .Y(_06851_),
    .A1(net624),
    .A2(_06850_));
 sg13g2_nor2_1 _12879_ (.A(net624),
    .B(_06850_),
    .Y(_06852_));
 sg13g2_or2_1 _12880_ (.X(_06853_),
    .B(_06852_),
    .A(_03110_));
 sg13g2_nand2_1 _12881_ (.Y(_06854_),
    .A(_03029_),
    .B(_03048_));
 sg13g2_nand2b_1 _12882_ (.Y(_06855_),
    .B(_04427_),
    .A_N(_06854_));
 sg13g2_nand2_1 _12883_ (.Y(_06856_),
    .A(_03007_),
    .B(_05835_));
 sg13g2_and2_1 _12884_ (.A(_06854_),
    .B(_05198_),
    .X(_06857_));
 sg13g2_a221oi_1 _12885_ (.B2(_06856_),
    .C1(_06857_),
    .B1(_06855_),
    .A1(net624),
    .Y(_06858_),
    .A2(_06850_));
 sg13g2_a21o_1 _12886_ (.A2(_06853_),
    .A1(_06851_),
    .B1(_06858_),
    .X(_06859_));
 sg13g2_nand2b_1 _12887_ (.Y(_06860_),
    .B(net623),
    .A_N(_03110_));
 sg13g2_nand3_1 _12888_ (.B(_06859_),
    .C(_06860_),
    .A(_06849_),
    .Y(_06861_));
 sg13g2_and3_1 _12889_ (.X(_06862_),
    .A(_02820_),
    .B(_05128_),
    .C(_05162_));
 sg13g2_buf_2 fanout460 (.A(net461),
    .X(net460));
 sg13g2_nor2_1 _12891_ (.A(_02781_),
    .B(net354),
    .Y(_06864_));
 sg13g2_nand2_1 _12892_ (.Y(_06865_),
    .A(_02670_),
    .B(_05237_));
 sg13g2_nor2_1 _12893_ (.A(_02729_),
    .B(_05120_),
    .Y(_06866_));
 sg13g2_a22oi_1 _12894_ (.Y(_06867_),
    .B1(_06865_),
    .B2(_06866_),
    .A2(net354),
    .A1(_02781_));
 sg13g2_nand4_1 _12895_ (.B(_05095_),
    .C(_05104_),
    .A(_02729_),
    .Y(_06868_),
    .D(_05118_));
 sg13g2_a21oi_1 _12896_ (.A1(_02781_),
    .A2(net354),
    .Y(_06869_),
    .B1(_06868_));
 sg13g2_or4_1 _12897_ (.A(_06862_),
    .B(_06864_),
    .C(_06867_),
    .D(_06869_),
    .X(_06870_));
 sg13g2_nor2_1 _12898_ (.A(_04832_),
    .B(_04830_),
    .Y(_06871_));
 sg13g2_a21oi_1 _12899_ (.A1(_02946_),
    .A2(net618),
    .Y(_06872_),
    .B1(_06871_));
 sg13g2_nor2_1 _12900_ (.A(_02946_),
    .B(net618),
    .Y(_06873_));
 sg13g2_nor2_1 _12901_ (.A(_02917_),
    .B(_04928_),
    .Y(_06874_));
 sg13g2_a22oi_1 _12902_ (.Y(_06875_),
    .B1(net617),
    .B2(_02876_),
    .A2(_04928_),
    .A1(_02917_));
 sg13g2_or3_1 _12903_ (.A(_06873_),
    .B(_06874_),
    .C(_06875_),
    .X(_06876_));
 sg13g2_nor2_1 _12904_ (.A(_02974_),
    .B(_05177_),
    .Y(_06877_));
 sg13g2_a21oi_1 _12905_ (.A1(_06872_),
    .A2(_06876_),
    .Y(_06878_),
    .B1(_06877_));
 sg13g2_inv_1 _12906_ (.Y(_06879_),
    .A(_02820_));
 sg13g2_nand2_1 _12907_ (.Y(_06880_),
    .A(_06879_),
    .B(_05917_));
 sg13g2_nand3_1 _12908_ (.B(_06878_),
    .C(_06880_),
    .A(_06870_),
    .Y(_06881_));
 sg13g2_nand2_1 _12909_ (.Y(_06882_),
    .A(_04832_),
    .B(_04830_));
 sg13g2_nand2_1 _12910_ (.Y(_06883_),
    .A(_02917_),
    .B(_04928_));
 sg13g2_nand2_1 _12911_ (.Y(_06884_),
    .A(_02876_),
    .B(net617));
 sg13g2_a22oi_1 _12912_ (.Y(_06885_),
    .B1(_06874_),
    .B2(_06873_),
    .A2(_06884_),
    .A1(_06883_));
 sg13g2_nand2b_1 _12913_ (.Y(_06886_),
    .B(_06872_),
    .A_N(_06885_));
 sg13g2_a22oi_1 _12914_ (.Y(_06887_),
    .B1(net620),
    .B2(_04782_),
    .A2(_06836_),
    .A1(_04725_));
 sg13g2_o21ai_1 _12915_ (.B1(_06841_),
    .Y(_06888_),
    .A1(_06838_),
    .A2(_06887_));
 sg13g2_nor4_1 _12916_ (.A(_06841_),
    .B(_06844_),
    .C(_06838_),
    .D(_06887_),
    .Y(_06889_));
 sg13g2_a22oi_1 _12917_ (.Y(_06890_),
    .B1(_06889_),
    .B2(_06848_),
    .A2(_06888_),
    .A1(_06846_));
 sg13g2_a21oi_1 _12918_ (.A1(_06882_),
    .A2(_06886_),
    .Y(_06891_),
    .B1(_06890_));
 sg13g2_nand4_1 _12919_ (.B(_06861_),
    .C(_06881_),
    .A(_06835_),
    .Y(_06892_),
    .D(_06891_));
 sg13g2_nand2_1 _12920_ (.Y(_06893_),
    .A(net160),
    .B(net603));
 sg13g2_nand2_1 _12921_ (.Y(_06894_),
    .A(net159),
    .B(_05434_));
 sg13g2_nor2_1 _12922_ (.A(net160),
    .B(net603),
    .Y(_06895_));
 sg13g2_a221oi_1 _12923_ (.B2(_06894_),
    .C1(_06895_),
    .B1(_06893_),
    .A1(_03613_),
    .Y(_06896_),
    .A2(net599));
 sg13g2_nand2_1 _12924_ (.Y(_06897_),
    .A(net162),
    .B(net600));
 sg13g2_o21ai_1 _12925_ (.B1(_06897_),
    .Y(_06898_),
    .A1(_03613_),
    .A2(net599));
 sg13g2_nor2_1 _12926_ (.A(net162),
    .B(net601),
    .Y(_06899_));
 sg13g2_inv_1 _12927_ (.Y(_06900_),
    .A(_06899_));
 sg13g2_o21ai_1 _12928_ (.B1(_06900_),
    .Y(_06901_),
    .A1(_06896_),
    .A2(_06898_));
 sg13g2_a21o_1 _12929_ (.A2(net354),
    .A1(_02781_),
    .B1(_05917_),
    .X(_06902_));
 sg13g2_nand2b_1 _12930_ (.Y(_06903_),
    .B(net566),
    .A_N(_02729_));
 sg13g2_nand3_1 _12931_ (.B(net613),
    .C(_06868_),
    .A(_05032_),
    .Y(_06904_));
 sg13g2_a22oi_1 _12932_ (.Y(_06905_),
    .B1(net402),
    .B2(_06862_),
    .A2(_06904_),
    .A1(_06903_));
 sg13g2_a21oi_1 _12933_ (.A1(_06879_),
    .A2(_06902_),
    .Y(_06906_),
    .B1(_06905_));
 sg13g2_a21oi_1 _12934_ (.A1(_06903_),
    .A2(_06904_),
    .Y(_06907_),
    .B1(_06862_));
 sg13g2_nor2_1 _12935_ (.A(_05163_),
    .B(net402),
    .Y(_06908_));
 sg13g2_o21ai_1 _12936_ (.B1(_02781_),
    .Y(_06909_),
    .A1(_06907_),
    .A2(_06908_));
 sg13g2_nand4_1 _12937_ (.B(_06878_),
    .C(_06906_),
    .A(_06901_),
    .Y(_06910_),
    .D(_06909_));
 sg13g2_a22oi_1 _12938_ (.Y(_06911_),
    .B1(_05434_),
    .B2(net159),
    .A2(net603),
    .A1(net160));
 sg13g2_o21ai_1 _12939_ (.B1(net602),
    .Y(_06912_),
    .A1(net162),
    .A2(net600));
 sg13g2_nor3_1 _12940_ (.A(_06895_),
    .B(_06911_),
    .C(_06912_),
    .Y(_06913_));
 sg13g2_nor4_1 _12941_ (.A(_03613_),
    .B(_06899_),
    .C(_06895_),
    .D(_06911_),
    .Y(_06914_));
 sg13g2_o21ai_1 _12942_ (.B1(_06897_),
    .Y(_06915_),
    .A1(_03613_),
    .A2(_06912_));
 sg13g2_nor3_1 _12943_ (.A(_06913_),
    .B(_06914_),
    .C(_06915_),
    .Y(_06916_));
 sg13g2_nor2_1 _12944_ (.A(net144),
    .B(_05639_),
    .Y(_06917_));
 sg13g2_or2_1 _12945_ (.X(_06918_),
    .B(net648),
    .A(_03448_));
 sg13g2_nand2_1 _12946_ (.Y(_06919_),
    .A(net144),
    .B(_05639_));
 sg13g2_o21ai_1 _12947_ (.B1(_06919_),
    .Y(_06920_),
    .A1(_06917_),
    .A2(_06918_));
 sg13g2_inv_1 _12948_ (.Y(_06921_),
    .A(net144));
 sg13g2_or2_1 _12949_ (.X(_06922_),
    .B(_05656_),
    .A(_06921_));
 sg13g2_a22oi_1 _12950_ (.Y(_06923_),
    .B1(_03501_),
    .B2(_06917_),
    .A2(_06922_),
    .A1(_06918_));
 sg13g2_nand2_1 _12951_ (.Y(_06924_),
    .A(net155),
    .B(_05776_));
 sg13g2_o21ai_1 _12952_ (.B1(_06924_),
    .Y(_06925_),
    .A1(_03543_),
    .A2(net391));
 sg13g2_a22oi_1 _12953_ (.Y(_06926_),
    .B1(_06923_),
    .B2(_06925_),
    .A2(_06920_),
    .A1(_05776_));
 sg13g2_a22oi_1 _12954_ (.Y(_06927_),
    .B1(_06916_),
    .B2(_06926_),
    .A2(net391),
    .A1(_03543_));
 sg13g2_nor2_1 _12955_ (.A(_06910_),
    .B(_06927_),
    .Y(_06928_));
 sg13g2_nor2_1 _12956_ (.A(_03007_),
    .B(_05835_),
    .Y(_06929_));
 sg13g2_a221oi_1 _12957_ (.B2(_06929_),
    .C1(_06857_),
    .B1(_06855_),
    .A1(net624),
    .Y(_06930_),
    .A2(_06850_));
 sg13g2_o21ai_1 _12958_ (.B1(net612),
    .Y(_06931_),
    .A1(_06852_),
    .A2(_06930_));
 sg13g2_o21ai_1 _12959_ (.B1(_03110_),
    .Y(_06932_),
    .A1(_06851_),
    .A2(_06930_));
 sg13g2_nand3b_1 _12960_ (.B(_06931_),
    .C(_06932_),
    .Y(_06933_),
    .A_N(_06890_));
 sg13g2_nand2b_1 _12961_ (.Y(_06934_),
    .B(_03989_),
    .A_N(_03889_));
 sg13g2_inv_1 _12962_ (.Y(_06935_),
    .A(_06827_));
 sg13g2_nand2_1 _12963_ (.Y(_06936_),
    .A(_06824_),
    .B(net568));
 sg13g2_nor2b_1 _12964_ (.A(net632),
    .B_N(_03296_),
    .Y(_06937_));
 sg13g2_a21oi_1 _12965_ (.A1(_06823_),
    .A2(_06936_),
    .Y(_06938_),
    .B1(_06937_));
 sg13g2_o21ai_1 _12966_ (.B1(_06822_),
    .Y(_06939_),
    .A1(_06935_),
    .A2(_06938_));
 sg13g2_and4_1 _12967_ (.A(_06819_),
    .B(_06934_),
    .C(_06849_),
    .D(_06939_),
    .X(_06940_));
 sg13g2_a21o_1 _12968_ (.A2(_06830_),
    .A1(_06819_),
    .B1(_06834_),
    .X(_06941_));
 sg13g2_a21o_1 _12969_ (.A2(_06940_),
    .A1(_06933_),
    .B1(_06941_),
    .X(_06942_));
 sg13g2_o21ai_1 _12970_ (.B1(_06942_),
    .Y(_06943_),
    .A1(_06892_),
    .A2(_06928_));
 sg13g2_xor2_1 _12971_ (.B(_06943_),
    .A(net1242),
    .X(_06944_));
 sg13g2_and4_1 _12972_ (.A(net1248),
    .B(net1237),
    .C(_05446_),
    .D(_02570_),
    .X(_06945_));
 sg13g2_and2_1 _12973_ (.A(_06933_),
    .B(_06940_),
    .X(_06946_));
 sg13g2_and2_1 _12974_ (.A(_03448_),
    .B(net647),
    .X(_06947_));
 sg13g2_a21oi_1 _12975_ (.A1(_06919_),
    .A2(_06947_),
    .Y(_06948_),
    .B1(_06917_));
 sg13g2_nand2_1 _12976_ (.Y(_06949_),
    .A(_03543_),
    .B(net598));
 sg13g2_nor4_1 _12977_ (.A(net155),
    .B(_05534_),
    .C(_05545_),
    .D(_05561_),
    .Y(_06950_));
 sg13g2_o21ai_1 _12978_ (.B1(_06950_),
    .Y(_06951_),
    .A1(_03543_),
    .A2(net598));
 sg13g2_a21o_1 _12979_ (.A2(_06951_),
    .A1(_06949_),
    .B1(net895),
    .X(_06952_));
 sg13g2_o21ai_1 _12980_ (.B1(_06952_),
    .Y(_06953_),
    .A1(_06925_),
    .A2(_06948_));
 sg13g2_and2_1 _12981_ (.A(_06901_),
    .B(_06953_),
    .X(_06954_));
 sg13g2_nor4_1 _12982_ (.A(_06916_),
    .B(_06954_),
    .C(_06910_),
    .D(_06927_),
    .Y(_06955_));
 sg13g2_inv_1 _12983_ (.Y(_06956_),
    .A(_03816_));
 sg13g2_nor3_1 _12984_ (.A(net1237),
    .B(net1239),
    .C(_06956_),
    .Y(_06957_));
 sg13g2_and2_1 _12985_ (.A(net1242),
    .B(_06957_),
    .X(_06958_));
 sg13g2_inv_1 _12986_ (.Y(_06959_),
    .A(_06958_));
 sg13g2_a21oi_1 _12987_ (.A1(_06946_),
    .A2(_06955_),
    .Y(_06960_),
    .B1(_06959_));
 sg13g2_and4_1 _12988_ (.A(_06835_),
    .B(_06861_),
    .C(_06881_),
    .D(_06891_),
    .X(_06961_));
 sg13g2_nor2b_1 _12989_ (.A(net1242),
    .B_N(_06957_),
    .Y(_06962_));
 sg13g2_nand4_1 _12990_ (.B(_06946_),
    .C(_06955_),
    .A(_06961_),
    .Y(_06963_),
    .D(_06962_));
 sg13g2_a21oi_1 _12991_ (.A1(_06892_),
    .A2(_06958_),
    .Y(_06964_),
    .B1(_03826_));
 sg13g2_nand3b_1 _12992_ (.B(_06963_),
    .C(_06964_),
    .Y(_06965_),
    .A_N(_06960_));
 sg13g2_a21oi_1 _12993_ (.A1(_06944_),
    .A2(_06945_),
    .Y(_06966_),
    .B1(_06965_));
 sg13g2_buf_2 fanout459 (.A(net462),
    .X(net459));
 sg13g2_buf_1 fanout458 (.A(net459),
    .X(net458));
 sg13g2_buf_2 fanout457 (.A(net459),
    .X(net457));
 sg13g2_buf_1 fanout456 (.A(_02329_),
    .X(net456));
 sg13g2_mux2_1 _12998_ (.A0(_06804_),
    .A1(_01024_),
    .S(net335),
    .X(\dp.ISRmux.d0[2] ));
 sg13g2_buf_2 fanout455 (.A(net456),
    .X(net455));
 sg13g2_nor2_1 _13000_ (.A(_01025_),
    .B(net884),
    .Y(_06972_));
 sg13g2_a21oi_1 _13001_ (.A1(net598),
    .A2(_06780_),
    .Y(_06973_),
    .B1(_06972_));
 sg13g2_xnor2_1 _13002_ (.Y(_06974_),
    .A(net871),
    .B(_06973_));
 sg13g2_a21oi_1 _13003_ (.A1(_05591_),
    .A2(_06780_),
    .Y(_06975_),
    .B1(_06799_));
 sg13g2_a21o_1 _13004_ (.A2(_05505_),
    .A1(_05504_),
    .B1(_05510_),
    .X(_06976_));
 sg13g2_a21o_1 _13005_ (.A2(_06975_),
    .A1(_06794_),
    .B1(_06976_),
    .X(_06977_));
 sg13g2_o21ai_1 _13006_ (.B1(_06977_),
    .Y(_06978_),
    .A1(_06794_),
    .A2(_06975_));
 sg13g2_xor2_1 _13007_ (.B(_06978_),
    .A(_06974_),
    .X(_06979_));
 sg13g2_xor2_1 _13008_ (.B(net122),
    .A(net125),
    .X(_06980_));
 sg13g2_mux2_1 _13009_ (.A0(_06979_),
    .A1(_06980_),
    .S(net335),
    .X(\dp.ISRmux.d0[3] ));
 sg13g2_buf_2 fanout454 (.A(net455),
    .X(net454));
 sg13g2_buf_2 fanout453 (.A(net456),
    .X(net453));
 sg13g2_inv_1 _13012_ (.Y(_06983_),
    .A(_01025_));
 sg13g2_o21ai_1 _13013_ (.B1(_05567_),
    .Y(_06984_),
    .A1(_06983_),
    .A2(net871));
 sg13g2_nand2_1 _13014_ (.Y(_06985_),
    .A(_06983_),
    .B(net871));
 sg13g2_o21ai_1 _13015_ (.B1(_06985_),
    .Y(_06986_),
    .A1(_01024_),
    .A2(_06984_));
 sg13g2_nor4_1 _13016_ (.A(_06785_),
    .B(_06793_),
    .C(_06801_),
    .D(_06802_),
    .Y(_06987_));
 sg13g2_nand2_1 _13017_ (.Y(_06988_),
    .A(net598),
    .B(_06780_));
 sg13g2_a21oi_1 _13018_ (.A1(_01024_),
    .A2(net892),
    .Y(_06989_),
    .B1(_06976_));
 sg13g2_nand3_1 _13019_ (.B(_05563_),
    .C(_06989_),
    .A(net871),
    .Y(_06990_));
 sg13g2_a21oi_1 _13020_ (.A1(_05563_),
    .A2(_06989_),
    .Y(_06991_),
    .B1(_05453_));
 sg13g2_a21oi_1 _13021_ (.A1(_06988_),
    .A2(_06990_),
    .Y(_06992_),
    .B1(_06991_));
 sg13g2_a221oi_1 _13022_ (.B2(_06974_),
    .C1(_06992_),
    .B1(_06987_),
    .A1(net892),
    .Y(_06993_),
    .A2(_06986_));
 sg13g2_buf_2 fanout452 (.A(net456),
    .X(net452));
 sg13g2_nor2_1 _13024_ (.A(_01026_),
    .B(net885),
    .Y(_06995_));
 sg13g2_a21oi_1 _13025_ (.A1(_05276_),
    .A2(net885),
    .Y(_06996_),
    .B1(_06995_));
 sg13g2_xnor2_1 _13026_ (.Y(_06997_),
    .A(_05876_),
    .B(_06996_));
 sg13g2_xor2_1 _13027_ (.B(_06997_),
    .A(_06993_),
    .X(_06998_));
 sg13g2_nand2_1 _13028_ (.Y(_06999_),
    .A(net125),
    .B(net122));
 sg13g2_xnor2_1 _13029_ (.Y(_07000_),
    .A(net126),
    .B(_06999_));
 sg13g2_mux2_1 _13030_ (.A0(_06998_),
    .A1(_07000_),
    .S(net333),
    .X(\dp.ISRmux.d0[4] ));
 sg13g2_nand2_1 _13031_ (.Y(_07001_),
    .A(_01027_),
    .B(net893));
 sg13g2_o21ai_1 _13032_ (.B1(_07001_),
    .Y(_07002_),
    .A1(_06076_),
    .A2(net893));
 sg13g2_xnor2_1 _13033_ (.Y(_07003_),
    .A(_05319_),
    .B(_07002_));
 sg13g2_a21o_1 _13034_ (.A2(_06993_),
    .A1(_05876_),
    .B1(_06996_),
    .X(_07004_));
 sg13g2_o21ai_1 _13035_ (.B1(_07004_),
    .Y(_07005_),
    .A1(_05876_),
    .A2(_06993_));
 sg13g2_xnor2_1 _13036_ (.Y(_07006_),
    .A(_07003_),
    .B(_07005_));
 sg13g2_nor2_1 _13037_ (.A(_01026_),
    .B(_06999_),
    .Y(_07007_));
 sg13g2_xor2_1 _13038_ (.B(_07007_),
    .A(net127),
    .X(_07008_));
 sg13g2_mux2_1 _13039_ (.A0(_07006_),
    .A1(_07008_),
    .S(net333),
    .X(\dp.ISRmux.d0[5] ));
 sg13g2_nor2_1 _13040_ (.A(_05876_),
    .B(net892),
    .Y(_07009_));
 sg13g2_nor2b_1 _13041_ (.A(_05876_),
    .B_N(_06995_),
    .Y(_07010_));
 sg13g2_a221oi_1 _13042_ (.B2(_07009_),
    .C1(_07010_),
    .B1(_05276_),
    .A1(net18),
    .Y(_07011_),
    .A2(net942));
 sg13g2_inv_1 _13043_ (.Y(_07012_),
    .A(_01026_));
 sg13g2_nor2_1 _13044_ (.A(_05876_),
    .B(_05319_),
    .Y(_07013_));
 sg13g2_a21oi_1 _13045_ (.A1(_07012_),
    .A2(_07013_),
    .Y(_07014_),
    .B1(_07001_));
 sg13g2_a22oi_1 _13046_ (.Y(_07015_),
    .B1(net893),
    .B2(_06076_),
    .A2(_07013_),
    .A1(_05276_));
 sg13g2_nor3_1 _13047_ (.A(_07011_),
    .B(_07014_),
    .C(_07015_),
    .Y(_07016_));
 sg13g2_or3_1 _13048_ (.A(_06993_),
    .B(_06997_),
    .C(_07003_),
    .X(_07017_));
 sg13g2_nand2b_1 _13049_ (.Y(_07018_),
    .B(_07017_),
    .A_N(_07016_));
 sg13g2_buf_2 fanout451 (.A(net456),
    .X(net451));
 sg13g2_and2_1 _13051_ (.A(_01028_),
    .B(net892),
    .X(_07020_));
 sg13g2_a22oi_1 _13052_ (.Y(_07021_),
    .B1(_07020_),
    .B2(_05368_),
    .A2(net885),
    .A1(net602));
 sg13g2_nor2_1 _13053_ (.A(_01028_),
    .B(net885),
    .Y(_07022_));
 sg13g2_a22oi_1 _13054_ (.Y(_07023_),
    .B1(_07022_),
    .B2(_05364_),
    .A2(net885),
    .A1(net599));
 sg13g2_or2_1 _13055_ (.X(_07024_),
    .B(_07023_),
    .A(_07021_));
 sg13g2_xnor2_1 _13056_ (.Y(_07025_),
    .A(_07018_),
    .B(_07024_));
 sg13g2_nand4_1 _13057_ (.B(net122),
    .C(net126),
    .A(net125),
    .Y(_07026_),
    .D(net127));
 sg13g2_buf_2 fanout450 (.A(net451),
    .X(net450));
 sg13g2_xnor2_1 _13059_ (.Y(_07028_),
    .A(net128),
    .B(_07026_));
 sg13g2_mux2_1 _13060_ (.A0(_07025_),
    .A1(_07028_),
    .S(net333),
    .X(\dp.ISRmux.d0[6] ));
 sg13g2_and2_1 _13061_ (.A(_01029_),
    .B(net892),
    .X(_07029_));
 sg13g2_a22oi_1 _13062_ (.Y(_07030_),
    .B1(_07029_),
    .B2(_05328_),
    .A2(net884),
    .A1(net601));
 sg13g2_o21ai_1 _13063_ (.B1(_05328_),
    .Y(_07031_),
    .A1(_01029_),
    .A2(net884));
 sg13g2_a21oi_1 _13064_ (.A1(_05362_),
    .A2(net884),
    .Y(_07032_),
    .B1(_07031_));
 sg13g2_or2_1 _13065_ (.X(_07033_),
    .B(_07032_),
    .A(_07030_));
 sg13g2_buf_2 fanout449 (.A(net451),
    .X(net449));
 sg13g2_a21oi_1 _13067_ (.A1(net599),
    .A2(net885),
    .Y(_07035_),
    .B1(_07022_));
 sg13g2_nor2_1 _13068_ (.A(_05364_),
    .B(_07018_),
    .Y(_07036_));
 sg13g2_nand2_1 _13069_ (.Y(_07037_),
    .A(_05364_),
    .B(_07018_));
 sg13g2_o21ai_1 _13070_ (.B1(_07037_),
    .Y(_07038_),
    .A1(_07035_),
    .A2(_07036_));
 sg13g2_xnor2_1 _13071_ (.Y(_07039_),
    .A(_07033_),
    .B(_07038_));
 sg13g2_nor2_1 _13072_ (.A(_01028_),
    .B(_07026_),
    .Y(_07040_));
 sg13g2_xor2_1 _13073_ (.B(_07040_),
    .A(net129),
    .X(_07041_));
 sg13g2_mux2_1 _13074_ (.A0(_07039_),
    .A1(_07041_),
    .S(net333),
    .X(\dp.ISRmux.d0[7] ));
 sg13g2_or4_1 _13075_ (.A(_06997_),
    .B(_07003_),
    .C(_07024_),
    .D(_07033_),
    .X(_07042_));
 sg13g2_nor4_1 _13076_ (.A(_07021_),
    .B(_07023_),
    .C(_07030_),
    .D(_07032_),
    .Y(_07043_));
 sg13g2_nor3_1 _13077_ (.A(_05368_),
    .B(_07035_),
    .C(_07032_),
    .Y(_07044_));
 sg13g2_a22oi_1 _13078_ (.Y(_07045_),
    .B1(_07044_),
    .B2(_07030_),
    .A2(_07043_),
    .A1(_07016_));
 sg13g2_o21ai_1 _13079_ (.B1(_07045_),
    .Y(_07046_),
    .A1(_06993_),
    .A2(_07042_));
 sg13g2_buf_2 fanout448 (.A(net449),
    .X(net448));
 sg13g2_nor2_1 _13081_ (.A(_01030_),
    .B(net886),
    .Y(_07048_));
 sg13g2_a21oi_1 _13082_ (.A1(_05237_),
    .A2(net886),
    .Y(_07049_),
    .B1(_07048_));
 sg13g2_xnor2_1 _13083_ (.Y(_07050_),
    .A(_05028_),
    .B(_07049_));
 sg13g2_xnor2_1 _13084_ (.Y(_07051_),
    .A(_07046_),
    .B(_07050_));
 sg13g2_nand2_1 _13085_ (.Y(_07052_),
    .A(net128),
    .B(net129));
 sg13g2_or2_1 _13086_ (.X(_07053_),
    .B(_07052_),
    .A(_07026_));
 sg13g2_buf_2 fanout447 (.A(net449),
    .X(net447));
 sg13g2_xnor2_1 _13088_ (.Y(_07055_),
    .A(net130),
    .B(_07053_));
 sg13g2_mux2_1 _13089_ (.A0(_07051_),
    .A1(_07055_),
    .S(net336),
    .X(\dp.ISRmux.d0[8] ));
 sg13g2_nand2_1 _13090_ (.Y(_07056_),
    .A(_01031_),
    .B(net893));
 sg13g2_o21ai_1 _13091_ (.B1(_07056_),
    .Y(_07057_),
    .A1(_05120_),
    .A2(net893));
 sg13g2_xnor2_1 _13092_ (.Y(_07058_),
    .A(_04987_),
    .B(_07057_));
 sg13g2_nor2b_1 _13093_ (.A(_07046_),
    .B_N(_05028_),
    .Y(_07059_));
 sg13g2_nand2b_1 _13094_ (.Y(_07060_),
    .B(_07046_),
    .A_N(_05028_));
 sg13g2_o21ai_1 _13095_ (.B1(_07060_),
    .Y(_07061_),
    .A1(_07049_),
    .A2(_07059_));
 sg13g2_xnor2_1 _13096_ (.Y(_07062_),
    .A(_07058_),
    .B(_07061_));
 sg13g2_nor2_1 _13097_ (.A(_01030_),
    .B(_07053_),
    .Y(_07063_));
 sg13g2_xor2_1 _13098_ (.B(_07063_),
    .A(net131),
    .X(_07064_));
 sg13g2_buf_1 fanout446 (.A(_02367_),
    .X(net446));
 sg13g2_mux2_1 _13100_ (.A0(_07062_),
    .A1(_07064_),
    .S(net336),
    .X(\dp.ISRmux.d0[9] ));
 sg13g2_or2_1 _13101_ (.X(_07066_),
    .B(_07058_),
    .A(_07050_));
 sg13g2_buf_1 fanout445 (.A(net446),
    .X(net445));
 sg13g2_inv_1 _13103_ (.Y(_07068_),
    .A(_07066_));
 sg13g2_nand2b_1 _13104_ (.Y(_07069_),
    .B(net21),
    .A_N(_01030_));
 sg13g2_nor2_1 _13105_ (.A(_01031_),
    .B(_07069_),
    .Y(_07070_));
 sg13g2_nor2_1 _13106_ (.A(net22),
    .B(_07070_),
    .Y(_07071_));
 sg13g2_a21oi_1 _13107_ (.A1(_01031_),
    .A2(_07069_),
    .Y(_07072_),
    .B1(_07071_));
 sg13g2_o21ai_1 _13108_ (.B1(net940),
    .Y(_07073_),
    .A1(_05449_),
    .A2(_07072_));
 sg13g2_nand2_1 _13109_ (.Y(_07074_),
    .A(net567),
    .B(net886));
 sg13g2_o21ai_1 _13110_ (.B1(_04186_),
    .Y(_07075_),
    .A1(net886),
    .A2(_07069_));
 sg13g2_and2_1 _13111_ (.A(_04987_),
    .B(net886),
    .X(_07076_));
 sg13g2_a22oi_1 _13112_ (.Y(_07077_),
    .B1(_04280_),
    .B2(net614),
    .A2(_07076_),
    .A1(net567));
 sg13g2_a21oi_1 _13113_ (.A1(_07074_),
    .A2(_07075_),
    .Y(_07078_),
    .B1(_07077_));
 sg13g2_nor2_1 _13114_ (.A(_07073_),
    .B(_07078_),
    .Y(_07079_));
 sg13g2_a21oi_1 _13115_ (.A1(_07046_),
    .A2(_07068_),
    .Y(_07080_),
    .B1(_07079_));
 sg13g2_a21oi_1 _13116_ (.A1(net942),
    .A2(_05082_),
    .Y(_07081_),
    .B1(_06789_));
 sg13g2_nor2_1 _13117_ (.A(_01032_),
    .B(net884),
    .Y(_07082_));
 sg13g2_a21o_2 _13118_ (.A2(_07081_),
    .A1(_05058_),
    .B1(_07082_),
    .X(_07083_));
 sg13g2_buf_2 fanout444 (.A(net445),
    .X(net444));
 sg13g2_xor2_1 _13120_ (.B(_07083_),
    .A(_04982_),
    .X(_07085_));
 sg13g2_xnor2_1 _13121_ (.Y(_07086_),
    .A(_07080_),
    .B(_07085_));
 sg13g2_inv_1 _13122_ (.Y(_07087_),
    .A(_07053_));
 sg13g2_nand3_1 _13123_ (.B(net131),
    .C(_07087_),
    .A(net130),
    .Y(_07088_));
 sg13g2_buf_2 fanout443 (.A(net446),
    .X(net443));
 sg13g2_xnor2_1 _13125_ (.Y(_07090_),
    .A(net101),
    .B(_07088_));
 sg13g2_mux2_1 _13126_ (.A0(_07086_),
    .A1(_07090_),
    .S(net334),
    .X(\dp.ISRmux.d0[10] ));
 sg13g2_and2_1 _13127_ (.A(_05128_),
    .B(net884),
    .X(_07091_));
 sg13g2_nor2_1 _13128_ (.A(_01033_),
    .B(net884),
    .Y(_07092_));
 sg13g2_mux2_1 _13129_ (.A0(_07092_),
    .A1(_01033_),
    .S(_05167_),
    .X(_07093_));
 sg13g2_a22oi_1 _13130_ (.Y(_07094_),
    .B1(_07093_),
    .B2(_05168_),
    .A2(_07091_),
    .A1(_05162_));
 sg13g2_a21o_1 _13131_ (.A2(_05168_),
    .A1(net401),
    .B1(_07094_),
    .X(_07095_));
 sg13g2_buf_2 fanout442 (.A(net446),
    .X(net442));
 sg13g2_a21o_1 _13133_ (.A2(_07068_),
    .A1(_07046_),
    .B1(_07079_),
    .X(_07097_));
 sg13g2_nor2_1 _13134_ (.A(_07097_),
    .B(_07083_),
    .Y(_07098_));
 sg13g2_a21oi_1 _13135_ (.A1(_07097_),
    .A2(_07083_),
    .Y(_07099_),
    .B1(_04982_));
 sg13g2_nor2_1 _13136_ (.A(_07098_),
    .B(_07099_),
    .Y(_07100_));
 sg13g2_xnor2_1 _13137_ (.Y(_07101_),
    .A(_07095_),
    .B(_07100_));
 sg13g2_nor2_1 _13138_ (.A(_01032_),
    .B(_07088_),
    .Y(_07102_));
 sg13g2_xor2_1 _13139_ (.B(_07102_),
    .A(net102),
    .X(_07103_));
 sg13g2_mux2_1 _13140_ (.A0(_07101_),
    .A1(_07103_),
    .S(net334),
    .X(\dp.ISRmux.d0[11] ));
 sg13g2_nand2b_1 _13141_ (.Y(_07104_),
    .B(_07085_),
    .A_N(_07095_));
 sg13g2_nor2_1 _13142_ (.A(_05167_),
    .B(_05168_),
    .Y(_07105_));
 sg13g2_nand2_1 _13143_ (.Y(_07106_),
    .A(_04982_),
    .B(_07083_));
 sg13g2_buf_1 fanout441 (.A(net446),
    .X(net441));
 sg13g2_nor2b_1 _13145_ (.A(_07105_),
    .B_N(_04982_),
    .Y(_07108_));
 sg13g2_a221oi_1 _13146_ (.B2(_07108_),
    .C1(_07092_),
    .B1(_07083_),
    .A1(net401),
    .Y(_07109_),
    .A2(net884));
 sg13g2_a21o_1 _13147_ (.A2(_07106_),
    .A1(_07105_),
    .B1(_07109_),
    .X(_07110_));
 sg13g2_buf_2 fanout440 (.A(net441),
    .X(net440));
 sg13g2_o21ai_1 _13149_ (.B1(_07110_),
    .Y(_07112_),
    .A1(_07080_),
    .A2(_07104_));
 sg13g2_buf_1 fanout439 (.A(net440),
    .X(net439));
 sg13g2_a21o_1 _13151_ (.A2(_04488_),
    .A1(net1243),
    .B1(net898),
    .X(_07114_));
 sg13g2_buf_2 fanout438 (.A(net440),
    .X(net438));
 sg13g2_nor2_1 _13153_ (.A(_01034_),
    .B(net887),
    .Y(_07116_));
 sg13g2_a21o_1 _13154_ (.A2(net887),
    .A1(net616),
    .B1(_07116_),
    .X(_07117_));
 sg13g2_buf_2 fanout437 (.A(net441),
    .X(net437));
 sg13g2_xnor2_1 _13156_ (.Y(_07119_),
    .A(_07114_),
    .B(_07117_));
 sg13g2_xnor2_1 _13157_ (.Y(_07120_),
    .A(_07112_),
    .B(_07119_));
 sg13g2_nand2_1 _13158_ (.Y(_07121_),
    .A(net101),
    .B(net102));
 sg13g2_nor2_1 _13159_ (.A(_07088_),
    .B(_07121_),
    .Y(_07122_));
 sg13g2_xor2_1 _13160_ (.B(_07122_),
    .A(net103),
    .X(_07123_));
 sg13g2_mux2_1 _13161_ (.A0(_07120_),
    .A1(_07123_),
    .S(net331),
    .X(\dp.ISRmux.d0[12] ));
 sg13g2_a21oi_1 _13162_ (.A1(net1241),
    .A2(net896),
    .Y(_07124_),
    .B1(net898));
 sg13g2_nand2b_1 _13163_ (.Y(_07125_),
    .B(net894),
    .A_N(_01035_));
 sg13g2_o21ai_1 _13164_ (.B1(_07125_),
    .Y(_07126_),
    .A1(_05185_),
    .A2(net894));
 sg13g2_xor2_1 _13165_ (.B(_07126_),
    .A(_07124_),
    .X(_07127_));
 sg13g2_a21o_1 _13166_ (.A2(_07117_),
    .A1(_07112_),
    .B1(_07114_),
    .X(_07128_));
 sg13g2_o21ai_1 _13167_ (.B1(_07128_),
    .Y(_07129_),
    .A1(_07112_),
    .A2(_07117_));
 sg13g2_xnor2_1 _13168_ (.Y(_07130_),
    .A(_07127_),
    .B(_07129_));
 sg13g2_nor3_1 _13169_ (.A(_01034_),
    .B(_07088_),
    .C(_07121_),
    .Y(_07131_));
 sg13g2_xor2_1 _13170_ (.B(_07131_),
    .A(net104),
    .X(_07132_));
 sg13g2_nand2_1 _13171_ (.Y(_07133_),
    .A(net331),
    .B(_07132_));
 sg13g2_o21ai_1 _13172_ (.B1(_07133_),
    .Y(\dp.ISRmux.d0[13] ),
    .A1(net331),
    .A2(_07130_));
 sg13g2_or2_1 _13173_ (.X(_07134_),
    .B(_07127_),
    .A(_07119_));
 sg13g2_buf_1 fanout436 (.A(net437),
    .X(net436));
 sg13g2_nor3_1 _13175_ (.A(_07066_),
    .B(_07104_),
    .C(_07134_),
    .Y(_07136_));
 sg13g2_nand3b_1 _13176_ (.B(_07114_),
    .C(_07116_),
    .Y(_07137_),
    .A_N(_01035_));
 sg13g2_a21oi_1 _13177_ (.A1(_07114_),
    .A2(_07117_),
    .Y(_07138_),
    .B1(_07126_));
 sg13g2_a21oi_1 _13178_ (.A1(_07124_),
    .A2(_07137_),
    .Y(_07139_),
    .B1(_07138_));
 sg13g2_xnor2_1 _13179_ (.Y(_07140_),
    .A(_04982_),
    .B(_07083_));
 sg13g2_or4_1 _13180_ (.A(_07073_),
    .B(_07078_),
    .C(_07140_),
    .D(_07095_),
    .X(_07141_));
 sg13g2_a21oi_1 _13181_ (.A1(_07110_),
    .A2(_07141_),
    .Y(_07142_),
    .B1(_07134_));
 sg13g2_a22oi_1 _13182_ (.Y(_07143_),
    .B1(_07139_),
    .B2(_07142_),
    .A2(_07136_),
    .A1(_07046_));
 sg13g2_buf_2 fanout435 (.A(net437),
    .X(net435));
 sg13g2_a21o_1 _13184_ (.A2(net896),
    .A1(net1238),
    .B1(net898),
    .X(_07145_));
 sg13g2_nor2_1 _13185_ (.A(_01036_),
    .B(net887),
    .Y(_07146_));
 sg13g2_a21oi_1 _13186_ (.A1(net619),
    .A2(net887),
    .Y(_07147_),
    .B1(_07146_));
 sg13g2_xnor2_1 _13187_ (.Y(_07148_),
    .A(_07145_),
    .B(_07147_));
 sg13g2_xnor2_1 _13188_ (.Y(_07149_),
    .A(_07143_),
    .B(_07148_));
 sg13g2_nand4_1 _13189_ (.B(net131),
    .C(net103),
    .A(net130),
    .Y(_07150_),
    .D(net104));
 sg13g2_nor3_2 _13190_ (.A(_07053_),
    .B(_07121_),
    .C(_07150_),
    .Y(_07151_));
 sg13g2_xor2_1 _13191_ (.B(_07151_),
    .A(net105),
    .X(_07152_));
 sg13g2_mux2_1 _13192_ (.A0(_07149_),
    .A1(_07152_),
    .S(net331),
    .X(\dp.ISRmux.d0[14] ));
 sg13g2_a22oi_1 _13193_ (.Y(_07153_),
    .B1(_04826_),
    .B2(_06789_),
    .A2(_04819_),
    .A1(_04815_));
 sg13g2_nand2_1 _13194_ (.Y(_07154_),
    .A(_04809_),
    .B(_07153_));
 sg13g2_o21ai_1 _13195_ (.B1(_07154_),
    .Y(_07155_),
    .A1(_01037_),
    .A2(net887));
 sg13g2_xor2_1 _13196_ (.B(_07155_),
    .A(_04834_),
    .X(_07156_));
 sg13g2_a21o_1 _13197_ (.A2(_07143_),
    .A1(_04839_),
    .B1(_07147_),
    .X(_07157_));
 sg13g2_o21ai_1 _13198_ (.B1(_07157_),
    .Y(_07158_),
    .A1(_04839_),
    .A2(_07143_));
 sg13g2_xor2_1 _13199_ (.B(_07158_),
    .A(_07156_),
    .X(_07159_));
 sg13g2_nor2b_1 _13200_ (.A(_01036_),
    .B_N(_07151_),
    .Y(_07160_));
 sg13g2_xor2_1 _13201_ (.B(_07160_),
    .A(net106),
    .X(_07161_));
 sg13g2_mux2_1 _13202_ (.A0(_07159_),
    .A1(_07161_),
    .S(net332),
    .X(\dp.ISRmux.d0[15] ));
 sg13g2_nand2b_1 _13203_ (.Y(_07162_),
    .B(net894),
    .A_N(_01038_));
 sg13g2_nand4_1 _13204_ (.B(_04528_),
    .C(_04548_),
    .A(_04517_),
    .Y(_07163_),
    .D(net887));
 sg13g2_and2_1 _13205_ (.A(_07162_),
    .B(_07163_),
    .X(_07164_));
 sg13g2_xnor2_1 _13206_ (.Y(_07165_),
    .A(_04505_),
    .B(_07164_));
 sg13g2_nand2_1 _13207_ (.Y(_07166_),
    .A(_07148_),
    .B(_07156_));
 sg13g2_nor4_1 _13208_ (.A(_07066_),
    .B(_07104_),
    .C(_07134_),
    .D(_07166_),
    .Y(_07167_));
 sg13g2_a21o_1 _13209_ (.A2(_07137_),
    .A1(_07124_),
    .B1(_07138_),
    .X(_07168_));
 sg13g2_nand2_1 _13210_ (.Y(_07169_),
    .A(net619),
    .B(net887));
 sg13g2_inv_1 _13211_ (.Y(_07170_),
    .A(_01037_));
 sg13g2_o21ai_1 _13212_ (.B1(_07146_),
    .Y(_07171_),
    .A1(_07170_),
    .A2(_04834_));
 sg13g2_a21oi_1 _13213_ (.A1(_07169_),
    .A2(_07171_),
    .Y(_07172_),
    .B1(_04839_));
 sg13g2_a21oi_1 _13214_ (.A1(_04834_),
    .A2(_07155_),
    .Y(_07173_),
    .B1(_07172_));
 sg13g2_o21ai_1 _13215_ (.B1(_07173_),
    .Y(_07174_),
    .A1(_07168_),
    .A2(_07166_));
 sg13g2_a22oi_1 _13216_ (.Y(_07175_),
    .B1(_07166_),
    .B2(_07134_),
    .A2(_07141_),
    .A1(_07110_));
 sg13g2_a22oi_1 _13217_ (.Y(_07176_),
    .B1(_07174_),
    .B2(_07175_),
    .A2(_07167_),
    .A1(_07046_));
 sg13g2_buf_1 fanout434 (.A(_02405_),
    .X(net434));
 sg13g2_xor2_1 _13219_ (.B(_07176_),
    .A(_07165_),
    .X(_07178_));
 sg13g2_nand3_1 _13220_ (.B(net106),
    .C(_07151_),
    .A(net105),
    .Y(_07179_));
 sg13g2_buf_2 fanout433 (.A(_02405_),
    .X(net433));
 sg13g2_xnor2_1 _13222_ (.Y(_07181_),
    .A(net107),
    .B(_07179_));
 sg13g2_mux2_1 _13223_ (.A0(_07178_),
    .A1(_07181_),
    .S(net331),
    .X(\dp.ISRmux.d0[16] ));
 sg13g2_a21oi_1 _13224_ (.A1(_07162_),
    .A2(_07163_),
    .Y(_07182_),
    .B1(_04505_));
 sg13g2_nor2_1 _13225_ (.A(_07165_),
    .B(_07176_),
    .Y(_07183_));
 sg13g2_nor2_1 _13226_ (.A(_07182_),
    .B(_07183_),
    .Y(_07184_));
 sg13g2_and2_1 _13227_ (.A(_01039_),
    .B(net891),
    .X(_07185_));
 sg13g2_nor2_1 _13228_ (.A(net897),
    .B(_04439_),
    .Y(_07186_));
 sg13g2_a22oi_1 _13229_ (.Y(_07187_),
    .B1(_07185_),
    .B2(_07186_),
    .A2(net888),
    .A1(_05198_));
 sg13g2_buf_2 fanout432 (.A(_02408_),
    .X(net432));
 sg13g2_nor3_1 _13231_ (.A(net897),
    .B(_04439_),
    .C(net891),
    .Y(_07189_));
 sg13g2_and2_1 _13232_ (.A(_07186_),
    .B(_07185_),
    .X(_07190_));
 sg13g2_a21oi_1 _13233_ (.A1(_05198_),
    .A2(_07189_),
    .Y(_07191_),
    .B1(_07190_));
 sg13g2_nand2b_1 _13234_ (.Y(_07192_),
    .B(_07191_),
    .A_N(_07187_));
 sg13g2_xor2_1 _13235_ (.B(_07192_),
    .A(_07184_),
    .X(_07193_));
 sg13g2_nor2_1 _13236_ (.A(_01038_),
    .B(_07179_),
    .Y(_07194_));
 sg13g2_xor2_1 _13237_ (.B(_07194_),
    .A(net108),
    .X(_07195_));
 sg13g2_mux2_1 _13238_ (.A0(_07193_),
    .A1(_07195_),
    .S(net329),
    .X(\dp.ISRmux.d0[17] ));
 sg13g2_and2_1 _13239_ (.A(_01040_),
    .B(net891),
    .X(_07196_));
 sg13g2_a21o_1 _13240_ (.A2(net883),
    .A1(net625),
    .B1(_07196_),
    .X(_07197_));
 sg13g2_xnor2_1 _13241_ (.Y(_07198_),
    .A(_04490_),
    .B(_07197_));
 sg13g2_nand2b_1 _13242_ (.Y(_07199_),
    .B(_07191_),
    .A_N(_07165_));
 sg13g2_o21ai_1 _13243_ (.B1(_07191_),
    .Y(_07200_),
    .A1(_07182_),
    .A2(_07187_));
 sg13g2_o21ai_1 _13244_ (.B1(_07200_),
    .Y(_07201_),
    .A1(_07176_),
    .A2(_07199_));
 sg13g2_buf_2 fanout431 (.A(net432),
    .X(net431));
 sg13g2_xnor2_1 _13246_ (.Y(_07203_),
    .A(_07198_),
    .B(_07201_));
 sg13g2_nand2_1 _13247_ (.Y(_07204_),
    .A(net107),
    .B(net108));
 sg13g2_or2_1 _13248_ (.X(_07205_),
    .B(_07204_),
    .A(_07179_));
 sg13g2_buf_2 fanout430 (.A(_02408_),
    .X(net430));
 sg13g2_xnor2_1 _13250_ (.Y(_07207_),
    .A(net109),
    .B(_07205_));
 sg13g2_mux2_1 _13251_ (.A0(_07203_),
    .A1(_07207_),
    .S(net329),
    .X(\dp.ISRmux.d0[18] ));
 sg13g2_a21oi_2 _13252_ (.B1(net897),
    .Y(_07208_),
    .A2(net896),
    .A1(net1395));
 sg13g2_nor2_1 _13253_ (.A(_01041_),
    .B(net883),
    .Y(_07209_));
 sg13g2_a21oi_1 _13254_ (.A1(net612),
    .A2(net888),
    .Y(_07210_),
    .B1(_07209_));
 sg13g2_xnor2_1 _13255_ (.Y(_07211_),
    .A(_07208_),
    .B(_07210_));
 sg13g2_inv_1 _13256_ (.Y(_07212_),
    .A(_07197_));
 sg13g2_nor2_1 _13257_ (.A(_07212_),
    .B(_07201_),
    .Y(_07213_));
 sg13g2_nand2_1 _13258_ (.Y(_07214_),
    .A(_07212_),
    .B(_07201_));
 sg13g2_o21ai_1 _13259_ (.B1(_07214_),
    .Y(_07215_),
    .A1(_04490_),
    .A2(_07213_));
 sg13g2_xnor2_1 _13260_ (.Y(_07216_),
    .A(_07211_),
    .B(_07215_));
 sg13g2_nor2_1 _13261_ (.A(_01040_),
    .B(_07205_),
    .Y(_07217_));
 sg13g2_xor2_1 _13262_ (.B(_07217_),
    .A(net110),
    .X(_07218_));
 sg13g2_mux2_1 _13263_ (.A0(_07216_),
    .A1(_07218_),
    .S(net329),
    .X(\dp.ISRmux.d0[19] ));
 sg13g2_or4_1 _13264_ (.A(_07165_),
    .B(_07192_),
    .C(_07198_),
    .D(_07211_),
    .X(_07219_));
 sg13g2_nor3_1 _13265_ (.A(_07198_),
    .B(_07200_),
    .C(_07211_),
    .Y(_07220_));
 sg13g2_or2_1 _13266_ (.X(_07221_),
    .B(_07196_),
    .A(_04490_));
 sg13g2_buf_2 fanout429 (.A(net430),
    .X(net429));
 sg13g2_nor2_1 _13268_ (.A(net625),
    .B(_07221_),
    .Y(_07223_));
 sg13g2_a21oi_1 _13269_ (.A1(net612),
    .A2(net888),
    .Y(_07224_),
    .B1(_07223_));
 sg13g2_a21oi_1 _13270_ (.A1(_07208_),
    .A2(_07221_),
    .Y(_07225_),
    .B1(_01041_));
 sg13g2_nor2_1 _13271_ (.A(_07208_),
    .B(_07221_),
    .Y(_07226_));
 sg13g2_o21ai_1 _13272_ (.B1(_06778_),
    .Y(_07227_),
    .A1(_07225_),
    .A2(_07226_));
 sg13g2_o21ai_1 _13273_ (.B1(_07227_),
    .Y(_07228_),
    .A1(_07208_),
    .A2(_07224_));
 sg13g2_nor2_1 _13274_ (.A(_07220_),
    .B(_07228_),
    .Y(_07229_));
 sg13g2_o21ai_1 _13275_ (.B1(_07229_),
    .Y(_07230_),
    .A1(_07176_),
    .A2(_07219_));
 sg13g2_buf_2 fanout428 (.A(_02408_),
    .X(net428));
 sg13g2_nor3_1 _13277_ (.A(_04758_),
    .B(_04778_),
    .C(net890),
    .Y(_07232_));
 sg13g2_a21oi_2 _13278_ (.B1(_07232_),
    .Y(_07233_),
    .A2(net890),
    .A1(_01042_));
 sg13g2_buf_2 fanout427 (.A(net428),
    .X(net427));
 sg13g2_xnor2_1 _13280_ (.Y(_07235_),
    .A(_04052_),
    .B(_07233_));
 sg13g2_xor2_1 _13281_ (.B(_07235_),
    .A(_07230_),
    .X(_07236_));
 sg13g2_nand2_1 _13282_ (.Y(_07237_),
    .A(net109),
    .B(net110));
 sg13g2_or2_1 _13283_ (.X(_07238_),
    .B(_07237_),
    .A(_07205_));
 sg13g2_buf_1 fanout426 (.A(net427),
    .X(net426));
 sg13g2_xnor2_1 _13285_ (.Y(_07240_),
    .A(net112),
    .B(_07238_));
 sg13g2_buf_2 fanout425 (.A(net427),
    .X(net425));
 sg13g2_mux2_1 _13287_ (.A0(_07236_),
    .A1(_07240_),
    .S(net325),
    .X(\dp.ISRmux.d0[20] ));
 sg13g2_a21oi_1 _13288_ (.A1(net1289),
    .A2(net918),
    .Y(_07242_),
    .B1(_03893_));
 sg13g2_and2_1 _13289_ (.A(_01043_),
    .B(net889),
    .X(_07243_));
 sg13g2_a21oi_2 _13290_ (.B1(_07243_),
    .Y(_07244_),
    .A2(net883),
    .A1(_04725_));
 sg13g2_xnor2_1 _13291_ (.Y(_07245_),
    .A(_07242_),
    .B(_07244_));
 sg13g2_a21o_1 _13292_ (.A2(_07233_),
    .A1(_07230_),
    .B1(_03895_),
    .X(_07246_));
 sg13g2_o21ai_1 _13293_ (.B1(_07246_),
    .Y(_07247_),
    .A1(_07230_),
    .A2(_07233_));
 sg13g2_xnor2_1 _13294_ (.Y(_07248_),
    .A(_07245_),
    .B(_07247_));
 sg13g2_nor2_1 _13295_ (.A(_01042_),
    .B(_07238_),
    .Y(_07249_));
 sg13g2_xor2_1 _13296_ (.B(_07249_),
    .A(net113),
    .X(_07250_));
 sg13g2_mux2_1 _13297_ (.A0(_07248_),
    .A1(_07250_),
    .S(net325),
    .X(\dp.ISRmux.d0[21] ));
 sg13g2_and2_1 _13298_ (.A(_01044_),
    .B(net889),
    .X(_07251_));
 sg13g2_a22oi_1 _13299_ (.Y(_07252_),
    .B1(_07251_),
    .B2(_04636_),
    .A2(net883),
    .A1(_05949_));
 sg13g2_nand2_1 _13300_ (.Y(_07253_),
    .A(_04636_),
    .B(net883));
 sg13g2_nand2_1 _13301_ (.Y(_07254_),
    .A(_04636_),
    .B(_07251_));
 sg13g2_o21ai_1 _13302_ (.B1(_07254_),
    .Y(_07255_),
    .A1(net622),
    .A2(_07253_));
 sg13g2_buf_1 fanout424 (.A(_02482_),
    .X(net424));
 sg13g2_nor2_1 _13304_ (.A(_07252_),
    .B(_07255_),
    .Y(_07257_));
 sg13g2_nor2_1 _13305_ (.A(_04729_),
    .B(_07244_),
    .Y(_07258_));
 sg13g2_a22oi_1 _13306_ (.Y(_07259_),
    .B1(_07233_),
    .B2(_03895_),
    .A2(_07244_),
    .A1(_04729_));
 sg13g2_nor2_1 _13307_ (.A(_07258_),
    .B(_07259_),
    .Y(_07260_));
 sg13g2_nand3_1 _13308_ (.B(_07233_),
    .C(_07244_),
    .A(_03895_),
    .Y(_07261_));
 sg13g2_a21oi_1 _13309_ (.A1(_03895_),
    .A2(_07233_),
    .Y(_07262_),
    .B1(_07244_));
 sg13g2_a21oi_1 _13310_ (.A1(_07242_),
    .A2(_07261_),
    .Y(_07263_),
    .B1(_07262_));
 sg13g2_a21oi_1 _13311_ (.A1(_07230_),
    .A2(_07260_),
    .Y(_07264_),
    .B1(_07263_));
 sg13g2_xnor2_1 _13312_ (.Y(_07265_),
    .A(_07257_),
    .B(_07264_));
 sg13g2_nand2_1 _13313_ (.Y(_07266_),
    .A(net112),
    .B(net113));
 sg13g2_nor2_1 _13314_ (.A(_07238_),
    .B(_07266_),
    .Y(_07267_));
 sg13g2_xor2_1 _13315_ (.B(_07267_),
    .A(net114),
    .X(_07268_));
 sg13g2_mux2_1 _13316_ (.A0(_07265_),
    .A1(_07268_),
    .S(net326),
    .X(\dp.ISRmux.d0[22] ));
 sg13g2_nand2_1 _13317_ (.Y(_07269_),
    .A(_01045_),
    .B(net889));
 sg13g2_o21ai_1 _13318_ (.B1(_07269_),
    .Y(_07270_),
    .A1(_04685_),
    .A2(net890));
 sg13g2_buf_1 fanout423 (.A(net424),
    .X(net423));
 sg13g2_xor2_1 _13320_ (.B(_07270_),
    .A(_04687_),
    .X(_07272_));
 sg13g2_a22oi_1 _13321_ (.Y(_07273_),
    .B1(_07263_),
    .B2(_07252_),
    .A2(_07260_),
    .A1(_07230_));
 sg13g2_or3_1 _13322_ (.A(_07255_),
    .B(_07272_),
    .C(_07273_),
    .X(_07274_));
 sg13g2_o21ai_1 _13323_ (.B1(_07272_),
    .Y(_07275_),
    .A1(_07255_),
    .A2(_07273_));
 sg13g2_nand2_1 _13324_ (.Y(_07276_),
    .A(_07274_),
    .B(_07275_));
 sg13g2_nor3_1 _13325_ (.A(_01044_),
    .B(_07238_),
    .C(_07266_),
    .Y(_07277_));
 sg13g2_xor2_1 _13326_ (.B(_07277_),
    .A(net115),
    .X(_07278_));
 sg13g2_mux2_1 _13327_ (.A0(_07276_),
    .A1(_07278_),
    .S(net325),
    .X(\dp.ISRmux.d0[23] ));
 sg13g2_and4_1 _13328_ (.A(_07235_),
    .B(_07245_),
    .C(_07257_),
    .D(_07272_),
    .X(_07279_));
 sg13g2_nand2b_1 _13329_ (.Y(_07280_),
    .B(_07279_),
    .A_N(_07219_));
 sg13g2_o21ai_1 _13330_ (.B1(_07279_),
    .Y(_07281_),
    .A1(_07220_),
    .A2(_07228_));
 sg13g2_a22oi_1 _13331_ (.Y(_07282_),
    .B1(_07262_),
    .B2(_07255_),
    .A2(_07261_),
    .A1(_07242_));
 sg13g2_nor2_1 _13332_ (.A(_04687_),
    .B(_07270_),
    .Y(_07283_));
 sg13g2_or2_1 _13333_ (.X(_07284_),
    .B(_07283_),
    .A(_07252_));
 sg13g2_nand2_1 _13334_ (.Y(_07285_),
    .A(_04687_),
    .B(_07270_));
 sg13g2_o21ai_1 _13335_ (.B1(_07285_),
    .Y(_07286_),
    .A1(_07282_),
    .A2(_07284_));
 sg13g2_and2_1 _13336_ (.A(_07281_),
    .B(_07286_),
    .X(_07287_));
 sg13g2_o21ai_1 _13337_ (.B1(_07287_),
    .Y(_07288_),
    .A1(_07176_),
    .A2(_07280_));
 sg13g2_buf_2 fanout422 (.A(net424),
    .X(net422));
 sg13g2_nand2_1 _13339_ (.Y(_07290_),
    .A(_05673_),
    .B(net883));
 sg13g2_nand2_1 _13340_ (.Y(_07291_),
    .A(_01046_),
    .B(net889));
 sg13g2_nand2_1 _13341_ (.Y(_07292_),
    .A(_07290_),
    .B(_07291_));
 sg13g2_xor2_1 _13342_ (.B(_07292_),
    .A(_04053_),
    .X(_07293_));
 sg13g2_xnor2_1 _13343_ (.Y(_07294_),
    .A(_07288_),
    .B(_07293_));
 sg13g2_and3_1 _13344_ (.X(_07295_),
    .A(net114),
    .B(net115),
    .C(_07267_));
 sg13g2_buf_2 fanout421 (.A(net424),
    .X(net421));
 sg13g2_xor2_1 _13346_ (.B(_07295_),
    .A(net116),
    .X(_07297_));
 sg13g2_mux2_1 _13347_ (.A0(_07294_),
    .A1(_07297_),
    .S(net326),
    .X(\dp.ISRmux.d0[24] ));
 sg13g2_nand2_1 _13348_ (.Y(_07298_),
    .A(net633),
    .B(net883));
 sg13g2_nand2_1 _13349_ (.Y(_07299_),
    .A(_01047_),
    .B(net889));
 sg13g2_a21oi_1 _13350_ (.A1(_07298_),
    .A2(_07299_),
    .Y(_07300_),
    .B1(_04106_));
 sg13g2_nand3_1 _13351_ (.B(_07298_),
    .C(_07299_),
    .A(_04106_),
    .Y(_07301_));
 sg13g2_buf_1 fanout420 (.A(net424),
    .X(net420));
 sg13g2_nand2b_1 _13353_ (.Y(_07303_),
    .B(_07301_),
    .A_N(_07300_));
 sg13g2_inv_1 _13354_ (.Y(_07304_),
    .A(_07292_));
 sg13g2_o21ai_1 _13355_ (.B1(_04053_),
    .Y(_07305_),
    .A1(_07288_),
    .A2(_07304_));
 sg13g2_nand2_1 _13356_ (.Y(_07306_),
    .A(_07288_),
    .B(_07304_));
 sg13g2_nand2_1 _13357_ (.Y(_07307_),
    .A(_07305_),
    .B(_07306_));
 sg13g2_xnor2_1 _13358_ (.Y(_07308_),
    .A(_07303_),
    .B(_07307_));
 sg13g2_nand2b_1 _13359_ (.Y(_07309_),
    .B(_07295_),
    .A_N(_01046_));
 sg13g2_xnor2_1 _13360_ (.Y(_07310_),
    .A(net117),
    .B(_07309_));
 sg13g2_mux2_1 _13361_ (.A0(_07308_),
    .A1(_07310_),
    .S(net326),
    .X(\dp.ISRmux.d0[25] ));
 sg13g2_nand3_1 _13362_ (.B(_07290_),
    .C(_07291_),
    .A(_04053_),
    .Y(_07311_));
 sg13g2_a21o_1 _13363_ (.A2(_07301_),
    .A1(_07311_),
    .B1(_07300_),
    .X(_07312_));
 sg13g2_or2_1 _13364_ (.X(_07313_),
    .B(_07303_),
    .A(_07293_));
 sg13g2_buf_2 fanout419 (.A(net420),
    .X(net419));
 sg13g2_nand2b_1 _13366_ (.Y(_07315_),
    .B(_07288_),
    .A_N(_07313_));
 sg13g2_nand2_1 _13367_ (.Y(_07316_),
    .A(_07312_),
    .B(_07315_));
 sg13g2_buf_2 fanout418 (.A(_02482_),
    .X(net418));
 sg13g2_nor2_1 _13369_ (.A(_05942_),
    .B(net890),
    .Y(_07318_));
 sg13g2_a21oi_2 _13370_ (.B1(_07318_),
    .Y(_07319_),
    .A2(net890),
    .A1(_01048_));
 sg13g2_xnor2_1 _13371_ (.Y(_07320_),
    .A(_04169_),
    .B(_07319_));
 sg13g2_xnor2_1 _13372_ (.Y(_07321_),
    .A(_07316_),
    .B(_07320_));
 sg13g2_and3_1 _13373_ (.X(_07322_),
    .A(net116),
    .B(net117),
    .C(_07295_));
 sg13g2_buf_2 fanout417 (.A(net418),
    .X(net417));
 sg13g2_xor2_1 _13375_ (.B(_07322_),
    .A(net118),
    .X(_07324_));
 sg13g2_mux2_1 _13376_ (.A0(_07321_),
    .A1(_07324_),
    .S(net327),
    .X(\dp.ISRmux.d0[26] ));
 sg13g2_and2_1 _13377_ (.A(_01049_),
    .B(net890),
    .X(_07325_));
 sg13g2_a21oi_1 _13378_ (.A1(_03989_),
    .A2(net883),
    .Y(_07326_),
    .B1(_07325_));
 sg13g2_nor2_1 _13379_ (.A(_03897_),
    .B(_07326_),
    .Y(_07327_));
 sg13g2_nand2_1 _13380_ (.Y(_07328_),
    .A(_03897_),
    .B(_07326_));
 sg13g2_nand2b_1 _13381_ (.Y(_07329_),
    .B(_07328_),
    .A_N(_07327_));
 sg13g2_a21oi_1 _13382_ (.A1(_07311_),
    .A2(_07301_),
    .Y(_07330_),
    .B1(_07300_));
 sg13g2_nor2_1 _13383_ (.A(_07330_),
    .B(_07319_),
    .Y(_07331_));
 sg13g2_nand3b_1 _13384_ (.B(_07312_),
    .C(_07313_),
    .Y(_07332_),
    .A_N(_04169_));
 sg13g2_o21ai_1 _13385_ (.B1(_07332_),
    .Y(_07333_),
    .A1(_04169_),
    .A2(_07319_));
 sg13g2_nor3_1 _13386_ (.A(_04169_),
    .B(_07288_),
    .C(_07330_),
    .Y(_07334_));
 sg13g2_a22oi_1 _13387_ (.Y(_07335_),
    .B1(_07333_),
    .B2(_07334_),
    .A2(_07331_),
    .A1(_07315_));
 sg13g2_xnor2_1 _13388_ (.Y(_07336_),
    .A(_07329_),
    .B(_07335_));
 sg13g2_nand2b_1 _13389_ (.Y(_07337_),
    .B(_07322_),
    .A_N(_01048_));
 sg13g2_xnor2_1 _13390_ (.Y(_07338_),
    .A(net119),
    .B(_07337_));
 sg13g2_mux2_1 _13391_ (.A0(_07336_),
    .A1(_07338_),
    .S(net327),
    .X(\dp.ISRmux.d0[27] ));
 sg13g2_nand2_1 _13392_ (.Y(_07339_),
    .A(_01050_),
    .B(net889));
 sg13g2_o21ai_1 _13393_ (.B1(_07339_),
    .Y(_07340_),
    .A1(_04278_),
    .A2(net891));
 sg13g2_xor2_1 _13394_ (.B(_07340_),
    .A(_04281_),
    .X(_07341_));
 sg13g2_or2_1 _13395_ (.X(_07342_),
    .B(_07329_),
    .A(_07320_));
 sg13g2_nor2_1 _13396_ (.A(_07313_),
    .B(_07342_),
    .Y(_07343_));
 sg13g2_a221oi_1 _13397_ (.B2(_03897_),
    .C1(_04169_),
    .B1(_07326_),
    .A1(_07330_),
    .Y(_07344_),
    .A2(_07319_));
 sg13g2_a22oi_1 _13398_ (.Y(_07345_),
    .B1(_07344_),
    .B2(_07327_),
    .A2(_07331_),
    .A1(_07328_));
 sg13g2_a21oi_1 _13399_ (.A1(_07288_),
    .A2(_07343_),
    .Y(_07346_),
    .B1(_07345_));
 sg13g2_xor2_1 _13400_ (.B(_07346_),
    .A(_07341_),
    .X(_07347_));
 sg13g2_nand3_1 _13401_ (.B(net119),
    .C(_07322_),
    .A(net118),
    .Y(_07348_));
 sg13g2_buf_2 fanout416 (.A(net418),
    .X(net416));
 sg13g2_xnor2_1 _13403_ (.Y(_07350_),
    .A(net120),
    .B(_07348_));
 sg13g2_mux2_1 _13404_ (.A0(_07347_),
    .A1(_07350_),
    .S(net328),
    .X(\dp.ISRmux.d0[28] ));
 sg13g2_nand2_1 _13405_ (.Y(_07351_),
    .A(_01051_),
    .B(net889));
 sg13g2_o21ai_1 _13406_ (.B1(_07351_),
    .Y(_07352_),
    .A1(_05868_),
    .A2(net889));
 sg13g2_buf_1 fanout415 (.A(net418),
    .X(net415));
 sg13g2_xor2_1 _13408_ (.B(_07352_),
    .A(_04187_),
    .X(_07354_));
 sg13g2_nor2b_1 _13409_ (.A(_07340_),
    .B_N(_04281_),
    .Y(_07355_));
 sg13g2_inv_1 _13410_ (.Y(_07356_),
    .A(_07355_));
 sg13g2_o21ai_1 _13411_ (.B1(_07356_),
    .Y(_07357_),
    .A1(_07341_),
    .A2(_07346_));
 sg13g2_xor2_1 _13412_ (.B(_07357_),
    .A(_07354_),
    .X(_07358_));
 sg13g2_nor2_1 _13413_ (.A(_01050_),
    .B(_07348_),
    .Y(_07359_));
 sg13g2_xor2_1 _13414_ (.B(_07359_),
    .A(net121),
    .X(_07360_));
 sg13g2_nand2_1 _13415_ (.Y(_07361_),
    .A(net328),
    .B(_07360_));
 sg13g2_o21ai_1 _13416_ (.B1(_07361_),
    .Y(\dp.ISRmux.d0[29] ),
    .A1(net328),
    .A2(_07358_));
 sg13g2_nor4_1 _13417_ (.A(_07313_),
    .B(_07341_),
    .C(_07342_),
    .D(_07354_),
    .Y(_07362_));
 sg13g2_nor2_1 _13418_ (.A(_07341_),
    .B(_07354_),
    .Y(_07363_));
 sg13g2_and2_1 _13419_ (.A(_07345_),
    .B(_07363_),
    .X(_07364_));
 sg13g2_nand2_1 _13420_ (.Y(_07365_),
    .A(_07356_),
    .B(_07352_));
 sg13g2_nor2_1 _13421_ (.A(_07356_),
    .B(_07352_),
    .Y(_07366_));
 sg13g2_a21oi_1 _13422_ (.A1(_04187_),
    .A2(_07365_),
    .Y(_07367_),
    .B1(_07366_));
 sg13g2_inv_1 _13423_ (.Y(_07368_),
    .A(_07367_));
 sg13g2_a22oi_1 _13424_ (.Y(_07369_),
    .B1(_07364_),
    .B2(_07368_),
    .A2(_07362_),
    .A1(_07288_));
 sg13g2_nor2_1 _13425_ (.A(_05684_),
    .B(net891),
    .Y(_07370_));
 sg13g2_a21oi_1 _13426_ (.A1(_01052_),
    .A2(net890),
    .Y(_07371_),
    .B1(_07370_));
 sg13g2_xnor2_1 _13427_ (.Y(_07372_),
    .A(_04392_),
    .B(_07371_));
 sg13g2_xor2_1 _13428_ (.B(_07372_),
    .A(_07369_),
    .X(_07373_));
 sg13g2_nand2_1 _13429_ (.Y(_07374_),
    .A(net120),
    .B(net121));
 sg13g2_nor2_1 _13430_ (.A(_07348_),
    .B(_07374_),
    .Y(_07375_));
 sg13g2_xor2_1 _13431_ (.B(_07375_),
    .A(net123),
    .X(_07376_));
 sg13g2_mux2_1 _13432_ (.A0(_07373_),
    .A1(_07376_),
    .S(net329),
    .X(\dp.ISRmux.d0[30] ));
 sg13g2_inv_1 _13433_ (.Y(_07377_),
    .A(_07371_));
 sg13g2_nor2_1 _13434_ (.A(_04392_),
    .B(_07371_),
    .Y(_07378_));
 sg13g2_nand2b_1 _13435_ (.Y(_07379_),
    .B(_07367_),
    .A_N(_04392_));
 sg13g2_a22oi_1 _13436_ (.Y(_07380_),
    .B1(_07364_),
    .B2(_07379_),
    .A2(_07362_),
    .A1(_07288_));
 sg13g2_a22oi_1 _13437_ (.Y(_07381_),
    .B1(_07378_),
    .B2(_07380_),
    .A2(_07377_),
    .A1(_07369_));
 sg13g2_nand2_1 _13438_ (.Y(_07382_),
    .A(net124),
    .B(net891));
 sg13g2_o21ai_1 _13439_ (.B1(_07382_),
    .Y(_07383_),
    .A1(net629),
    .A2(net891));
 sg13g2_xor2_1 _13440_ (.B(_07383_),
    .A(net25),
    .X(_07384_));
 sg13g2_xnor2_1 _13441_ (.Y(_07385_),
    .A(_07381_),
    .B(_07384_));
 sg13g2_nand2b_1 _13442_ (.Y(_07386_),
    .B(_07375_),
    .A_N(_01052_));
 sg13g2_xnor2_1 _13443_ (.Y(_07387_),
    .A(net124),
    .B(_07386_));
 sg13g2_nand2_1 _13444_ (.Y(_07388_),
    .A(net329),
    .B(_07387_));
 sg13g2_o21ai_1 _13445_ (.B1(_07388_),
    .Y(\dp.ISRmux.d0[31] ),
    .A1(net329),
    .A2(_07385_));
 sg13g2_nor4_1 _13446_ (.A(_02559_),
    .B(_03829_),
    .C(net986),
    .D(_03806_),
    .Y(net132));
 sg13g2_inv_1 _13447_ (.Y(_01053_),
    .A(net65));
 sg13g2_nor2_1 _13448_ (.A(net1256),
    .B(net1244),
    .Y(_07389_));
 sg13g2_and2_2 _13449_ (.A(net1247),
    .B(_07389_),
    .X(_07390_));
 sg13g2_buf_2 fanout414 (.A(net418),
    .X(net414));
 sg13g2_buf_1 fanout413 (.A(_02520_),
    .X(net413));
 sg13g2_a22oi_1 _13452_ (.Y(_07393_),
    .B1(_03826_),
    .B2(net919),
    .A2(_03870_),
    .A1(net985));
 sg13g2_buf_2 fanout412 (.A(net413),
    .X(net412));
 sg13g2_nor2_2 _13454_ (.A(_05645_),
    .B(_07393_),
    .Y(_07395_));
 sg13g2_and2_1 _13455_ (.A(net1245),
    .B(_07395_),
    .X(_07396_));
 sg13g2_buf_2 fanout411 (.A(_02520_),
    .X(net411));
 sg13g2_nand2_1 _13457_ (.Y(_07398_),
    .A(_07390_),
    .B(_07396_));
 sg13g2_buf_1 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_2 fanout409 (.A(net411),
    .X(net409));
 sg13g2_nor4_1 _13460_ (.A(net1252),
    .B(_03796_),
    .C(net1250),
    .D(net29),
    .Y(_07401_));
 sg13g2_a21o_1 _13461_ (.A2(_02561_),
    .A1(net29),
    .B1(_07401_),
    .X(_07402_));
 sg13g2_and3_1 _13462_ (.X(_07403_),
    .A(net1255),
    .B(_02565_),
    .C(_07402_));
 sg13g2_buf_2 fanout408 (.A(net411),
    .X(net408));
 sg13g2_nor2_1 _13464_ (.A(net828),
    .B(net861),
    .Y(_07405_));
 sg13g2_nor3_1 _13465_ (.A(net647),
    .B(_06786_),
    .C(net892),
    .Y(_07406_));
 sg13g2_and2_1 _13466_ (.A(net647),
    .B(_06786_),
    .X(_07407_));
 sg13g2_a22oi_1 _13467_ (.Y(_07408_),
    .B1(_07406_),
    .B2(_07407_),
    .A2(net892),
    .A1(_01022_));
 sg13g2_mux2_1 _13468_ (.A0(net100),
    .A1(_07408_),
    .S(net335),
    .X(_07409_));
 sg13g2_and2_1 _13469_ (.A(net860),
    .B(_07409_),
    .X(_07410_));
 sg13g2_a221oi_1 _13470_ (.B2(net66),
    .C1(_07410_),
    .B1(_07405_),
    .A1(net33),
    .Y(_07411_),
    .A2(net827));
 sg13g2_buf_2 fanout407 (.A(_02520_),
    .X(net407));
 sg13g2_buf_2 fanout406 (.A(net407),
    .X(net406));
 sg13g2_nand2_1 _13473_ (.Y(_07414_),
    .A(\dp.rf.rf[19][0] ),
    .B(net562));
 sg13g2_o21ai_1 _13474_ (.B1(_07414_),
    .Y(_01054_),
    .A1(net562),
    .A2(net302));
 sg13g2_buf_2 fanout405 (.A(net407),
    .X(net405));
 sg13g2_buf_2 fanout404 (.A(net407),
    .X(net404));
 sg13g2_buf_2 fanout403 (.A(_04977_),
    .X(net403));
 sg13g2_buf_2 fanout402 (.A(_05084_),
    .X(net402));
 sg13g2_buf_2 fanout401 (.A(_05163_),
    .X(net401));
 sg13g2_and2_1 _13480_ (.A(net44),
    .B(net827),
    .X(_07420_));
 sg13g2_a22oi_1 _13481_ (.Y(_07421_),
    .B1(net860),
    .B2(_07420_),
    .A2(net77),
    .A1(net867));
 sg13g2_a21oi_1 _13482_ (.A1(_05656_),
    .A2(_06780_),
    .Y(_07422_),
    .B1(_06783_));
 sg13g2_xnor2_1 _13483_ (.Y(_07423_),
    .A(_06788_),
    .B(_07407_));
 sg13g2_xnor2_1 _13484_ (.Y(_07424_),
    .A(_07422_),
    .B(_07423_));
 sg13g2_buf_2 fanout400 (.A(_05456_),
    .X(net400));
 sg13g2_nor2b_1 _13486_ (.A(net334),
    .B_N(net111),
    .Y(_07426_));
 sg13g2_nand3_1 _13487_ (.B(_02565_),
    .C(_07402_),
    .A(net1255),
    .Y(_07427_));
 sg13g2_buf_2 fanout399 (.A(net400),
    .X(net399));
 sg13g2_buf_1 fanout398 (.A(_05456_),
    .X(net398));
 sg13g2_a22oi_1 _13490_ (.Y(_07430_),
    .B1(_07426_),
    .B2(net855),
    .A2(_07424_),
    .A1(net334));
 sg13g2_or2_1 _13491_ (.X(_07431_),
    .B(_07430_),
    .A(_07421_));
 sg13g2_buf_2 fanout397 (.A(net398),
    .X(net397));
 sg13g2_buf_2 fanout396 (.A(net398),
    .X(net396));
 sg13g2_nand3_1 _13494_ (.B(_07390_),
    .C(_07395_),
    .A(net1245),
    .Y(_07434_));
 sg13g2_buf_2 fanout395 (.A(net396),
    .X(net395));
 sg13g2_buf_2 fanout394 (.A(_05456_),
    .X(net394));
 sg13g2_buf_1 fanout393 (.A(net394),
    .X(net393));
 sg13g2_nand2_1 _13498_ (.Y(_07438_),
    .A(\dp.rf.rf[19][1] ),
    .B(net812));
 sg13g2_o21ai_1 _13499_ (.B1(_07438_),
    .Y(_01055_),
    .A1(net297),
    .A2(net812));
 sg13g2_buf_2 fanout392 (.A(net394),
    .X(net392));
 sg13g2_buf_2 fanout391 (.A(_05498_),
    .X(net391));
 sg13g2_mux2_1 _13502_ (.A0(_01024_),
    .A1(_06804_),
    .S(net335),
    .X(_07441_));
 sg13g2_inv_1 _13503_ (.Y(_07442_),
    .A(net55));
 sg13g2_buf_1 fanout390 (.A(_05512_),
    .X(net390));
 sg13g2_nor2_1 _13505_ (.A(net827),
    .B(net88),
    .Y(_07444_));
 sg13g2_a22oi_1 _13506_ (.Y(_07445_),
    .B1(net860),
    .B2(_07444_),
    .A2(net827),
    .A1(_07442_));
 sg13g2_a21oi_1 _13507_ (.A1(net860),
    .A2(_07441_),
    .Y(_07446_),
    .B1(_07445_));
 sg13g2_buf_2 fanout389 (.A(net390),
    .X(net389));
 sg13g2_buf_1 fanout388 (.A(net390),
    .X(net388));
 sg13g2_nand2_1 _13510_ (.Y(_07449_),
    .A(\dp.rf.rf[19][2] ),
    .B(net813));
 sg13g2_o21ai_1 _13511_ (.B1(_07449_),
    .Y(_01056_),
    .A1(net812),
    .A2(net323));
 sg13g2_mux2_1 _13512_ (.A0(_06980_),
    .A1(_06979_),
    .S(net335),
    .X(_07450_));
 sg13g2_nand2_1 _13513_ (.Y(_07451_),
    .A(net58),
    .B(net827));
 sg13g2_nand2_1 _13514_ (.Y(_07452_),
    .A(net867),
    .B(net91));
 sg13g2_nand3_1 _13515_ (.B(_07451_),
    .C(_07452_),
    .A(net855),
    .Y(_07453_));
 sg13g2_o21ai_1 _13516_ (.B1(_07453_),
    .Y(_07454_),
    .A1(net856),
    .A2(_07450_));
 sg13g2_buf_2 fanout387 (.A(net388),
    .X(net387));
 sg13g2_buf_1 fanout386 (.A(_05512_),
    .X(net386));
 sg13g2_nand2_1 _13519_ (.Y(_07457_),
    .A(\dp.rf.rf[19][3] ),
    .B(net812));
 sg13g2_o21ai_1 _13520_ (.B1(_07457_),
    .Y(_01057_),
    .A1(net812),
    .A2(net318));
 sg13g2_mux2_1 _13521_ (.A0(_07000_),
    .A1(_06998_),
    .S(net333),
    .X(_07458_));
 sg13g2_inv_1 _13522_ (.Y(_07459_),
    .A(_07458_));
 sg13g2_and2_1 _13523_ (.A(net59),
    .B(net827),
    .X(_07460_));
 sg13g2_a22oi_1 _13524_ (.Y(_07461_),
    .B1(net859),
    .B2(_07460_),
    .A2(net92),
    .A1(net867));
 sg13g2_a21oi_1 _13525_ (.A1(net859),
    .A2(_07459_),
    .Y(_07462_),
    .B1(_07461_));
 sg13g2_buf_1 fanout385 (.A(net386),
    .X(net385));
 sg13g2_buf_2 fanout384 (.A(net385),
    .X(net384));
 sg13g2_mux2_1 _13528_ (.A0(net292),
    .A1(\dp.rf.rf[19][4] ),
    .S(net808),
    .X(_01058_));
 sg13g2_mux2_1 _13529_ (.A0(_07008_),
    .A1(_07006_),
    .S(net333),
    .X(_07465_));
 sg13g2_buf_2 fanout383 (.A(net385),
    .X(net383));
 sg13g2_and3_1 _13531_ (.X(_07467_),
    .A(net60),
    .B(net827),
    .C(net855));
 sg13g2_a221oi_1 _13532_ (.B2(net860),
    .C1(_07467_),
    .B1(_07465_),
    .A1(net93),
    .Y(_07468_),
    .A2(_07405_));
 sg13g2_buf_1 fanout382 (.A(net386),
    .X(net382));
 sg13g2_buf_2 fanout381 (.A(net386),
    .X(net381));
 sg13g2_nand2_1 _13535_ (.Y(_07471_),
    .A(\dp.rf.rf[19][5] ),
    .B(net810));
 sg13g2_o21ai_1 _13536_ (.B1(_07471_),
    .Y(_01059_),
    .A1(net810),
    .A2(net313));
 sg13g2_and2_1 _13537_ (.A(net61),
    .B(net828),
    .X(_07472_));
 sg13g2_a22oi_1 _13538_ (.Y(_07473_),
    .B1(net861),
    .B2(_07472_),
    .A2(net94),
    .A1(net866));
 sg13g2_mux2_1 _13539_ (.A0(_07028_),
    .A1(_07025_),
    .S(net333),
    .X(_07474_));
 sg13g2_nor2_1 _13540_ (.A(net855),
    .B(_07474_),
    .Y(_07475_));
 sg13g2_or2_1 _13541_ (.X(_07476_),
    .B(_07475_),
    .A(_07473_));
 sg13g2_buf_2 fanout380 (.A(net386),
    .X(net380));
 sg13g2_buf_2 fanout379 (.A(net380),
    .X(net379));
 sg13g2_nand2_1 _13544_ (.Y(_07479_),
    .A(\dp.rf.rf[19][6] ),
    .B(net810));
 sg13g2_o21ai_1 _13545_ (.B1(_07479_),
    .Y(_01060_),
    .A1(net810),
    .A2(net288));
 sg13g2_mux2_1 _13546_ (.A0(net62),
    .A1(net95),
    .S(net866),
    .X(_07480_));
 sg13g2_nand2_1 _13547_ (.Y(_07481_),
    .A(net334),
    .B(_07039_));
 sg13g2_nand2b_1 _13548_ (.Y(_07482_),
    .B(_07041_),
    .A_N(net333));
 sg13g2_a21oi_1 _13549_ (.A1(_07481_),
    .A2(_07482_),
    .Y(_07483_),
    .B1(net855));
 sg13g2_a21oi_2 _13550_ (.B1(_07483_),
    .Y(_07484_),
    .A2(_07480_),
    .A1(net855));
 sg13g2_buf_1 fanout378 (.A(_05516_),
    .X(net378));
 sg13g2_buf_1 fanout377 (.A(net378),
    .X(net377));
 sg13g2_nand2_1 _13553_ (.Y(_07487_),
    .A(\dp.rf.rf[19][7] ),
    .B(net811));
 sg13g2_o21ai_1 _13554_ (.B1(_07487_),
    .Y(_01061_),
    .A1(net811),
    .A2(net284));
 sg13g2_mux2_1 _13555_ (.A0(_07055_),
    .A1(_07051_),
    .S(net336),
    .X(_07488_));
 sg13g2_nand2_2 _13556_ (.Y(_07489_),
    .A(_02576_),
    .B(net828));
 sg13g2_buf_2 fanout376 (.A(net377),
    .X(net376));
 sg13g2_nand3b_1 _13558_ (.B(net62),
    .C(_02576_),
    .Y(_07491_),
    .A_N(net1238));
 sg13g2_nand2_1 _13559_ (.Y(_07492_),
    .A(net828),
    .B(_07491_));
 sg13g2_buf_2 fanout375 (.A(net376),
    .X(net375));
 sg13g2_a21oi_1 _13561_ (.A1(net63),
    .A2(_07489_),
    .Y(_07494_),
    .B1(net560));
 sg13g2_or2_1 _13562_ (.X(_07495_),
    .B(_07494_),
    .A(net859));
 sg13g2_a22oi_1 _13563_ (.Y(_07496_),
    .B1(_07495_),
    .B2(net833),
    .A2(_06188_),
    .A1(net867));
 sg13g2_nor2_1 _13564_ (.A(_06202_),
    .B(_07495_),
    .Y(_07497_));
 sg13g2_a22oi_1 _13565_ (.Y(_07498_),
    .B1(_07496_),
    .B2(_07497_),
    .A2(_07488_),
    .A1(net860));
 sg13g2_buf_2 fanout374 (.A(net378),
    .X(net374));
 sg13g2_buf_2 fanout373 (.A(net374),
    .X(net373));
 sg13g2_nand2_1 _13568_ (.Y(_07501_),
    .A(\dp.rf.rf[19][8] ),
    .B(net812));
 sg13g2_o21ai_1 _13569_ (.B1(_07501_),
    .Y(_01062_),
    .A1(net811),
    .A2(net279));
 sg13g2_mux2_1 _13570_ (.A0(_07064_),
    .A1(_07062_),
    .S(net336),
    .X(_07502_));
 sg13g2_buf_2 fanout372 (.A(net373),
    .X(net372));
 sg13g2_a21oi_1 _13572_ (.A1(net64),
    .A2(_07489_),
    .Y(_07504_),
    .B1(net561));
 sg13g2_or2_1 _13573_ (.X(_07505_),
    .B(_07504_),
    .A(_06217_));
 sg13g2_a22oi_1 _13574_ (.Y(_07506_),
    .B1(net859),
    .B2(_07505_),
    .A2(_06229_),
    .A1(net867));
 sg13g2_a21oi_2 _13575_ (.B1(_07506_),
    .Y(_07507_),
    .A2(_07502_),
    .A1(net859));
 sg13g2_buf_1 fanout371 (.A(net378),
    .X(net371));
 sg13g2_buf_2 fanout370 (.A(net371),
    .X(net370));
 sg13g2_nand2_1 _13578_ (.Y(_07510_),
    .A(\dp.rf.rf[19][9] ),
    .B(net562));
 sg13g2_o21ai_1 _13579_ (.B1(_07510_),
    .Y(_01063_),
    .A1(net562),
    .A2(net271));
 sg13g2_mux2_1 _13580_ (.A0(_07090_),
    .A1(_07086_),
    .S(net334),
    .X(_07511_));
 sg13g2_a22oi_1 _13581_ (.Y(_07512_),
    .B1(_06258_),
    .B2(net98),
    .A2(_06237_),
    .A1(net339));
 sg13g2_buf_2 fanout369 (.A(net371),
    .X(net369));
 sg13g2_a21oi_1 _13583_ (.A1(net34),
    .A2(_07489_),
    .Y(_07514_),
    .B1(net561));
 sg13g2_o21ai_1 _13584_ (.B1(net855),
    .Y(_07515_),
    .A1(_07512_),
    .A2(_07514_));
 sg13g2_o21ai_1 _13585_ (.B1(_07515_),
    .Y(_07516_),
    .A1(net856),
    .A2(_07511_));
 sg13g2_buf_1 fanout368 (.A(_05575_),
    .X(net368));
 sg13g2_buf_2 fanout367 (.A(net368),
    .X(net367));
 sg13g2_buf_2 fanout366 (.A(net367),
    .X(net366));
 sg13g2_nand2_1 _13589_ (.Y(_07520_),
    .A(\dp.rf.rf[19][10] ),
    .B(net810));
 sg13g2_o21ai_1 _13590_ (.B1(_07520_),
    .Y(_01064_),
    .A1(net810),
    .A2(net268));
 sg13g2_a21oi_1 _13591_ (.A1(net35),
    .A2(_07489_),
    .Y(_07521_),
    .B1(net560));
 sg13g2_nor2_1 _13592_ (.A(net859),
    .B(_07521_),
    .Y(_07522_));
 sg13g2_o21ai_1 _13593_ (.B1(_07522_),
    .Y(_07523_),
    .A1(net827),
    .A2(net68));
 sg13g2_mux2_1 _13594_ (.A0(_07103_),
    .A1(_07101_),
    .S(net334),
    .X(_07524_));
 sg13g2_nand2_1 _13595_ (.Y(_07525_),
    .A(net860),
    .B(_07524_));
 sg13g2_and2_1 _13596_ (.A(_07523_),
    .B(_07525_),
    .X(_07526_));
 sg13g2_buf_1 fanout365 (.A(net368),
    .X(net365));
 sg13g2_buf_2 fanout364 (.A(net365),
    .X(net364));
 sg13g2_nand2_1 _13599_ (.Y(_07529_),
    .A(\dp.rf.rf[19][11] ),
    .B(net812));
 sg13g2_o21ai_1 _13600_ (.B1(_07529_),
    .Y(_01065_),
    .A1(net812),
    .A2(net263));
 sg13g2_mux2_1 _13601_ (.A0(_07123_),
    .A1(_07120_),
    .S(net331),
    .X(_07530_));
 sg13g2_o21ai_1 _13602_ (.B1(net867),
    .Y(_07531_),
    .A1(_06296_),
    .A2(_06319_));
 sg13g2_a21o_1 _13603_ (.A2(_07489_),
    .A1(net36),
    .B1(net560),
    .X(_07532_));
 sg13g2_a21o_1 _13604_ (.A2(_07532_),
    .A1(_07531_),
    .B1(net859),
    .X(_07533_));
 sg13g2_o21ai_1 _13605_ (.B1(_07533_),
    .Y(_07534_),
    .A1(net855),
    .A2(_07530_));
 sg13g2_buf_1 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_2 fanout362 (.A(net364),
    .X(net362));
 sg13g2_nand2_1 _13608_ (.Y(_07537_),
    .A(\dp.rf.rf[19][12] ),
    .B(net810));
 sg13g2_o21ai_1 _13609_ (.B1(_07537_),
    .Y(_01066_),
    .A1(net810),
    .A2(net257));
 sg13g2_nand2b_1 _13610_ (.Y(_07538_),
    .B(net867),
    .A_N(net70));
 sg13g2_a21oi_1 _13611_ (.A1(net37),
    .A2(_07489_),
    .Y(_07539_),
    .B1(net561));
 sg13g2_nor2_1 _13612_ (.A(net859),
    .B(_07539_),
    .Y(_07540_));
 sg13g2_nor2_1 _13613_ (.A(net332),
    .B(_07132_),
    .Y(_07541_));
 sg13g2_a22oi_1 _13614_ (.Y(_07542_),
    .B1(_07541_),
    .B2(net856),
    .A2(_07130_),
    .A1(net332));
 sg13g2_a21o_1 _13615_ (.A2(_07540_),
    .A1(_07538_),
    .B1(_07542_),
    .X(_07543_));
 sg13g2_buf_2 fanout361 (.A(net365),
    .X(net361));
 sg13g2_buf_1 fanout360 (.A(net365),
    .X(net360));
 sg13g2_mux2_1 _13618_ (.A0(net250),
    .A1(\dp.rf.rf[19][13] ),
    .S(_07398_),
    .X(_01067_));
 sg13g2_mux2_1 _13619_ (.A0(_07152_),
    .A1(_07149_),
    .S(net331),
    .X(_07546_));
 sg13g2_a22oi_1 _13620_ (.Y(_07547_),
    .B1(_06370_),
    .B2(net828),
    .A2(_06348_),
    .A1(net339));
 sg13g2_a21oi_1 _13621_ (.A1(net38),
    .A2(_07489_),
    .Y(_07548_),
    .B1(net560));
 sg13g2_nor3_1 _13622_ (.A(net861),
    .B(_07547_),
    .C(_07548_),
    .Y(_07549_));
 sg13g2_a21oi_2 _13623_ (.B1(_07549_),
    .Y(_07550_),
    .A2(_07546_),
    .A1(net861));
 sg13g2_buf_2 fanout359 (.A(net360),
    .X(net359));
 sg13g2_buf_2 fanout358 (.A(_05788_),
    .X(net358));
 sg13g2_nand2_1 _13626_ (.Y(_07553_),
    .A(\dp.rf.rf[19][14] ),
    .B(net563));
 sg13g2_o21ai_1 _13627_ (.B1(_07553_),
    .Y(_01068_),
    .A1(net563),
    .A2(net246));
 sg13g2_mux2_1 _13628_ (.A0(_07161_),
    .A1(_07159_),
    .S(net332),
    .X(_07554_));
 sg13g2_nand3_1 _13629_ (.B(_06393_),
    .C(_07405_),
    .A(_06390_),
    .Y(_07555_));
 sg13g2_o21ai_1 _13630_ (.B1(_07555_),
    .Y(_07556_),
    .A1(net856),
    .A2(_07554_));
 sg13g2_a21oi_1 _13631_ (.A1(net39),
    .A2(_07489_),
    .Y(_07557_),
    .B1(net560));
 sg13g2_or2_1 _13632_ (.X(_07558_),
    .B(_07557_),
    .A(_07556_));
 sg13g2_buf_1 fanout357 (.A(_05800_),
    .X(net357));
 sg13g2_buf_2 fanout356 (.A(net357),
    .X(net356));
 sg13g2_nand2_1 _13635_ (.Y(_07561_),
    .A(\dp.rf.rf[19][15] ),
    .B(net562));
 sg13g2_o21ai_1 _13636_ (.B1(_07561_),
    .Y(_01069_),
    .A1(net562),
    .A2(net240));
 sg13g2_mux2_1 _13637_ (.A0(_07181_),
    .A1(_07178_),
    .S(net331),
    .X(_07562_));
 sg13g2_inv_1 _13638_ (.Y(_07563_),
    .A(net39));
 sg13g2_or4_1 _13639_ (.A(net6),
    .B(_07563_),
    .C(net983),
    .D(net866),
    .X(_07564_));
 sg13g2_buf_2 fanout355 (.A(net356),
    .X(net355));
 sg13g2_buf_2 fanout354 (.A(_05829_),
    .X(net354));
 sg13g2_buf_1 fanout353 (.A(_05879_),
    .X(net353));
 sg13g2_o21ai_1 _13643_ (.B1(net40),
    .Y(_07568_),
    .A1(net984),
    .A2(net866));
 sg13g2_and2_1 _13644_ (.A(_02576_),
    .B(net828),
    .X(_07569_));
 sg13g2_buf_1 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_1 fanout351 (.A(net352),
    .X(net351));
 sg13g2_a21oi_1 _13647_ (.A1(net805),
    .A2(_07568_),
    .Y(_07572_),
    .B1(net557));
 sg13g2_nor2_1 _13648_ (.A(net560),
    .B(_07572_),
    .Y(_07573_));
 sg13g2_nor2_1 _13649_ (.A(net828),
    .B(_06413_),
    .Y(_07574_));
 sg13g2_nor4_1 _13650_ (.A(_06403_),
    .B(net861),
    .C(_07573_),
    .D(_07574_),
    .Y(_07575_));
 sg13g2_a21oi_1 _13651_ (.A1(net861),
    .A2(_07562_),
    .Y(_07576_),
    .B1(_07575_));
 sg13g2_buf_2 fanout350 (.A(net352),
    .X(net350));
 sg13g2_buf_2 fanout349 (.A(net353),
    .X(net349));
 sg13g2_nand2_1 _13654_ (.Y(_07579_),
    .A(\dp.rf.rf[19][16] ),
    .B(net562));
 sg13g2_o21ai_1 _13655_ (.B1(_07579_),
    .Y(_01070_),
    .A1(net562),
    .A2(net234));
 sg13g2_buf_1 fanout348 (.A(net349),
    .X(net348));
 sg13g2_mux2_1 _13657_ (.A0(_07195_),
    .A1(_07193_),
    .S(net329),
    .X(_07581_));
 sg13g2_o21ai_1 _13658_ (.B1(net41),
    .Y(_07582_),
    .A1(net984),
    .A2(net866));
 sg13g2_a21oi_1 _13659_ (.A1(net805),
    .A2(_07582_),
    .Y(_07583_),
    .B1(net557));
 sg13g2_o21ai_1 _13660_ (.B1(net856),
    .Y(_07584_),
    .A1(net560),
    .A2(_07583_));
 sg13g2_a22oi_1 _13661_ (.Y(_07585_),
    .B1(_07584_),
    .B2(_06426_),
    .A2(_06435_),
    .A1(net866));
 sg13g2_a21oi_1 _13662_ (.A1(net861),
    .A2(_07581_),
    .Y(_07586_),
    .B1(_07585_));
 sg13g2_buf_2 fanout347 (.A(net349),
    .X(net347));
 sg13g2_buf_2 fanout346 (.A(_06022_),
    .X(net346));
 sg13g2_nand2_1 _13665_ (.Y(_07589_),
    .A(\dp.rf.rf[19][17] ),
    .B(net809));
 sg13g2_o21ai_1 _13666_ (.B1(_07589_),
    .Y(_01071_),
    .A1(net809),
    .A2(net232));
 sg13g2_o21ai_1 _13667_ (.B1(net42),
    .Y(_07590_),
    .A1(net983),
    .A2(net866));
 sg13g2_a21oi_1 _13668_ (.A1(net805),
    .A2(_07590_),
    .Y(_07591_),
    .B1(net557));
 sg13g2_nor2_1 _13669_ (.A(net560),
    .B(_07591_),
    .Y(_07592_));
 sg13g2_nor2_1 _13670_ (.A(net832),
    .B(_07592_),
    .Y(_07593_));
 sg13g2_a21o_1 _13671_ (.A2(_07593_),
    .A1(_06449_),
    .B1(_06458_),
    .X(_07594_));
 sg13g2_nor2_1 _13672_ (.A(net865),
    .B(_07592_),
    .Y(_07595_));
 sg13g2_nand2_1 _13673_ (.Y(_07596_),
    .A(net330),
    .B(_07203_));
 sg13g2_nand2b_1 _13674_ (.Y(_07597_),
    .B(_07207_),
    .A_N(net329));
 sg13g2_a21oi_1 _13675_ (.A1(_07596_),
    .A2(_07597_),
    .Y(_07598_),
    .B1(net854));
 sg13g2_a22oi_1 _13676_ (.Y(_07599_),
    .B1(_07595_),
    .B2(_07598_),
    .A2(_07594_),
    .A1(net854));
 sg13g2_buf_2 fanout345 (.A(net346),
    .X(net345));
 sg13g2_buf_2 fanout344 (.A(net345),
    .X(net344));
 sg13g2_nand2_1 _13679_ (.Y(_07602_),
    .A(\dp.rf.rf[19][18] ),
    .B(net811));
 sg13g2_o21ai_1 _13680_ (.B1(_07602_),
    .Y(_01072_),
    .A1(net811),
    .A2(net227));
 sg13g2_mux2_1 _13681_ (.A0(_07218_),
    .A1(_07216_),
    .S(net330),
    .X(_07603_));
 sg13g2_o21ai_1 _13682_ (.B1(net43),
    .Y(_07604_),
    .A1(net984),
    .A2(net866));
 sg13g2_a21oi_1 _13683_ (.A1(_07564_),
    .A2(_07604_),
    .Y(_07605_),
    .B1(_07569_));
 sg13g2_o21ai_1 _13684_ (.B1(net854),
    .Y(_07606_),
    .A1(net559),
    .A2(_07605_));
 sg13g2_a22oi_1 _13685_ (.Y(_07607_),
    .B1(_07606_),
    .B2(_06466_),
    .A2(_06479_),
    .A1(net865));
 sg13g2_a21oi_2 _13686_ (.B1(_07607_),
    .Y(_07608_),
    .A2(_07603_),
    .A1(net858));
 sg13g2_buf_2 fanout343 (.A(_06289_),
    .X(net343));
 sg13g2_buf_2 fanout342 (.A(_05793_),
    .X(net342));
 sg13g2_nand2_1 _13689_ (.Y(_07611_),
    .A(\dp.rf.rf[19][19] ),
    .B(net808));
 sg13g2_o21ai_1 _13690_ (.B1(_07611_),
    .Y(_01073_),
    .A1(net808),
    .A2(net222));
 sg13g2_a21o_1 _13691_ (.A2(_06504_),
    .A1(_06492_),
    .B1(net829),
    .X(_07612_));
 sg13g2_o21ai_1 _13692_ (.B1(net45),
    .Y(_07613_),
    .A1(net983),
    .A2(net864));
 sg13g2_a21oi_1 _13693_ (.A1(net804),
    .A2(_07613_),
    .Y(_07614_),
    .B1(net556));
 sg13g2_nor2_1 _13694_ (.A(net558),
    .B(_07614_),
    .Y(_07615_));
 sg13g2_nor2_1 _13695_ (.A(net857),
    .B(_07615_),
    .Y(_07616_));
 sg13g2_nor2b_1 _13696_ (.A(_07236_),
    .B_N(net325),
    .Y(_07617_));
 sg13g2_nor2_1 _13697_ (.A(net326),
    .B(_07240_),
    .Y(_07618_));
 sg13g2_nor3_1 _13698_ (.A(net853),
    .B(_07617_),
    .C(_07618_),
    .Y(_07619_));
 sg13g2_a21oi_1 _13699_ (.A1(_07612_),
    .A2(_07616_),
    .Y(_07620_),
    .B1(_07619_));
 sg13g2_buf_2 fanout341 (.A(_05818_),
    .X(net341));
 sg13g2_buf_2 fanout340 (.A(_06043_),
    .X(net340));
 sg13g2_nand2_1 _13702_ (.Y(_07623_),
    .A(\dp.rf.rf[19][20] ),
    .B(net806));
 sg13g2_o21ai_1 _13703_ (.B1(_07623_),
    .Y(_01074_),
    .A1(net806),
    .A2(net217));
 sg13g2_o21ai_1 _13704_ (.B1(net46),
    .Y(_07624_),
    .A1(net982),
    .A2(net864));
 sg13g2_a21oi_1 _13705_ (.A1(net805),
    .A2(_07624_),
    .Y(_07625_),
    .B1(net557));
 sg13g2_or2_1 _13706_ (.X(_07626_),
    .B(_07625_),
    .A(net559));
 sg13g2_o21ai_1 _13707_ (.B1(_07626_),
    .Y(_07627_),
    .A1(net829),
    .A2(net79));
 sg13g2_nor2b_1 _13708_ (.A(net325),
    .B_N(_07250_),
    .Y(_07628_));
 sg13g2_a21oi_1 _13709_ (.A1(net325),
    .A2(_07248_),
    .Y(_07629_),
    .B1(_07628_));
 sg13g2_mux2_1 _13710_ (.A0(_07627_),
    .A1(_07629_),
    .S(net857),
    .X(_07630_));
 sg13g2_buf_2 fanout339 (.A(_06141_),
    .X(net339));
 sg13g2_buf_2 fanout338 (.A(_05669_),
    .X(net338));
 sg13g2_nand2_1 _13713_ (.Y(_07633_),
    .A(\dp.rf.rf[19][21] ),
    .B(net806));
 sg13g2_o21ai_1 _13714_ (.B1(_07633_),
    .Y(_01075_),
    .A1(net806),
    .A2(net210));
 sg13g2_mux2_1 _13715_ (.A0(_07268_),
    .A1(_07265_),
    .S(net326),
    .X(_07634_));
 sg13g2_o21ai_1 _13716_ (.B1(net47),
    .Y(_07635_),
    .A1(net984),
    .A2(net865));
 sg13g2_a21oi_1 _13717_ (.A1(net805),
    .A2(_07635_),
    .Y(_07636_),
    .B1(net557));
 sg13g2_nor2_1 _13718_ (.A(net559),
    .B(_07636_),
    .Y(_07637_));
 sg13g2_a22oi_1 _13719_ (.Y(_07638_),
    .B1(net858),
    .B2(_07637_),
    .A2(_06559_),
    .A1(net865));
 sg13g2_a21oi_1 _13720_ (.A1(net857),
    .A2(_07634_),
    .Y(_07639_),
    .B1(_07638_));
 sg13g2_buf_1 fanout337 (.A(_06966_),
    .X(net337));
 sg13g2_buf_2 fanout336 (.A(net337),
    .X(net336));
 sg13g2_nand2_1 _13723_ (.Y(_07642_),
    .A(\dp.rf.rf[19][22] ),
    .B(net809));
 sg13g2_o21ai_1 _13724_ (.B1(_07642_),
    .Y(_01076_),
    .A1(net813),
    .A2(net208));
 sg13g2_and3_1 _13725_ (.X(_07643_),
    .A(net325),
    .B(_07274_),
    .C(_07275_));
 sg13g2_nor2_1 _13726_ (.A(net325),
    .B(_07278_),
    .Y(_07644_));
 sg13g2_nor3_1 _13727_ (.A(net853),
    .B(_07643_),
    .C(_07644_),
    .Y(_07645_));
 sg13g2_a21o_1 _13728_ (.A2(net854),
    .A1(net81),
    .B1(net829),
    .X(_07646_));
 sg13g2_o21ai_1 _13729_ (.B1(net48),
    .Y(_07647_),
    .A1(net983),
    .A2(net865));
 sg13g2_a21oi_1 _13730_ (.A1(net805),
    .A2(_07647_),
    .Y(_07648_),
    .B1(net557));
 sg13g2_or2_1 _13731_ (.X(_07649_),
    .B(_07648_),
    .A(net559));
 sg13g2_o21ai_1 _13732_ (.B1(_07649_),
    .Y(_07650_),
    .A1(_07645_),
    .A2(_07646_));
 sg13g2_buf_2 fanout335 (.A(net336),
    .X(net335));
 sg13g2_buf_2 fanout334 (.A(net335),
    .X(net334));
 sg13g2_nand2_1 _13735_ (.Y(_07653_),
    .A(\dp.rf.rf[19][23] ),
    .B(net563));
 sg13g2_o21ai_1 _13736_ (.B1(_07653_),
    .Y(_01077_),
    .A1(net563),
    .A2(net202));
 sg13g2_mux2_1 _13737_ (.A0(_07297_),
    .A1(_07294_),
    .S(net326),
    .X(_07654_));
 sg13g2_a22oi_1 _13738_ (.Y(_07655_),
    .B1(_06603_),
    .B2(net829),
    .A2(_06598_),
    .A1(net344));
 sg13g2_o21ai_1 _13739_ (.B1(net49),
    .Y(_07656_),
    .A1(net982),
    .A2(net862));
 sg13g2_a21oi_1 _13740_ (.A1(net804),
    .A2(_07656_),
    .Y(_07657_),
    .B1(net556));
 sg13g2_o21ai_1 _13741_ (.B1(net853),
    .Y(_07658_),
    .A1(net558),
    .A2(_07657_));
 sg13g2_nor3_1 _13742_ (.A(_06597_),
    .B(_07655_),
    .C(_07658_),
    .Y(_07659_));
 sg13g2_a21oi_1 _13743_ (.A1(net857),
    .A2(_07654_),
    .Y(_07660_),
    .B1(_07659_));
 sg13g2_buf_2 fanout333 (.A(net334),
    .X(net333));
 sg13g2_buf_1 fanout332 (.A(net337),
    .X(net332));
 sg13g2_nand2_1 _13746_ (.Y(_07663_),
    .A(\dp.rf.rf[19][24] ),
    .B(net807));
 sg13g2_o21ai_1 _13747_ (.B1(_07663_),
    .Y(_01078_),
    .A1(net807),
    .A2(net196));
 sg13g2_mux2_1 _13748_ (.A0(_07310_),
    .A1(_07308_),
    .S(net326),
    .X(_07664_));
 sg13g2_nor2_1 _13749_ (.A(_05671_),
    .B(net829),
    .Y(_07665_));
 sg13g2_and4_1 _13750_ (.A(_06605_),
    .B(_06607_),
    .C(_06630_),
    .D(_07665_),
    .X(_07666_));
 sg13g2_nand3_1 _13751_ (.B(net863),
    .C(_06630_),
    .A(_05671_),
    .Y(_07667_));
 sg13g2_nor2_1 _13752_ (.A(_06605_),
    .B(_07667_),
    .Y(_07668_));
 sg13g2_nand3_1 _13753_ (.B(net340),
    .C(_06630_),
    .A(net863),
    .Y(_07669_));
 sg13g2_o21ai_1 _13754_ (.B1(_07669_),
    .Y(_07670_),
    .A1(_06607_),
    .A2(_07667_));
 sg13g2_o21ai_1 _13755_ (.B1(net50),
    .Y(_07671_),
    .A1(net982),
    .A2(net862));
 sg13g2_a21oi_1 _13756_ (.A1(net804),
    .A2(_07671_),
    .Y(_07672_),
    .B1(net556));
 sg13g2_nor2_1 _13757_ (.A(net558),
    .B(_07672_),
    .Y(_07673_));
 sg13g2_nor2_1 _13758_ (.A(net857),
    .B(_07673_),
    .Y(_07674_));
 sg13g2_inv_1 _13759_ (.Y(_07675_),
    .A(_07674_));
 sg13g2_nor4_1 _13760_ (.A(_07666_),
    .B(_07668_),
    .C(_07670_),
    .D(_07675_),
    .Y(_07676_));
 sg13g2_a21oi_1 _13761_ (.A1(net857),
    .A2(_07664_),
    .Y(_07677_),
    .B1(_07676_));
 sg13g2_buf_2 fanout331 (.A(net337),
    .X(net331));
 sg13g2_buf_1 fanout330 (.A(net337),
    .X(net330));
 sg13g2_nand2_1 _13764_ (.Y(_07680_),
    .A(\dp.rf.rf[19][25] ),
    .B(net806));
 sg13g2_o21ai_1 _13765_ (.B1(_07680_),
    .Y(_01079_),
    .A1(net806),
    .A2(net191));
 sg13g2_mux2_1 _13766_ (.A0(_07324_),
    .A1(_07321_),
    .S(net327),
    .X(_07681_));
 sg13g2_o21ai_1 _13767_ (.B1(net51),
    .Y(_07682_),
    .A1(net982),
    .A2(net862));
 sg13g2_a21oi_1 _13768_ (.A1(net804),
    .A2(_07682_),
    .Y(_07683_),
    .B1(net556));
 sg13g2_nor2_1 _13769_ (.A(net558),
    .B(_07683_),
    .Y(_07684_));
 sg13g2_a22oi_1 _13770_ (.Y(_07685_),
    .B1(net857),
    .B2(_07684_),
    .A2(_06656_),
    .A1(net862));
 sg13g2_a21oi_1 _13771_ (.A1(net857),
    .A2(_07681_),
    .Y(_07686_),
    .B1(_07685_));
 sg13g2_buf_2 fanout329 (.A(net330),
    .X(net329));
 sg13g2_buf_2 fanout328 (.A(net330),
    .X(net328));
 sg13g2_nand2_1 _13774_ (.Y(_07689_),
    .A(\dp.rf.rf[19][26] ),
    .B(net563));
 sg13g2_o21ai_1 _13775_ (.B1(_07689_),
    .Y(_01080_),
    .A1(net563),
    .A2(net185));
 sg13g2_mux2_1 _13776_ (.A0(_07338_),
    .A1(_07336_),
    .S(net327),
    .X(_07690_));
 sg13g2_o21ai_1 _13777_ (.B1(net52),
    .Y(_07691_),
    .A1(net982),
    .A2(net862));
 sg13g2_a21oi_1 _13778_ (.A1(net804),
    .A2(_07691_),
    .Y(_07692_),
    .B1(net556));
 sg13g2_nor2_1 _13779_ (.A(net558),
    .B(_07692_),
    .Y(_07693_));
 sg13g2_nor2_1 _13780_ (.A(net863),
    .B(_07693_),
    .Y(_07694_));
 sg13g2_o21ai_1 _13781_ (.B1(net853),
    .Y(_07695_),
    .A1(net558),
    .A2(_07692_));
 sg13g2_a22oi_1 _13782_ (.Y(_07696_),
    .B1(_06681_),
    .B2(_07695_),
    .A2(_06669_),
    .A1(_06666_));
 sg13g2_a22oi_1 _13783_ (.Y(_07697_),
    .B1(_07694_),
    .B2(_07696_),
    .A2(_07690_),
    .A1(net858));
 sg13g2_buf_2 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_2 fanout326 (.A(net327),
    .X(net326));
 sg13g2_nand2_1 _13786_ (.Y(_07700_),
    .A(\dp.rf.rf[19][27] ),
    .B(net806));
 sg13g2_o21ai_1 _13787_ (.B1(_07700_),
    .Y(_01081_),
    .A1(net806),
    .A2(_07697_));
 sg13g2_mux2_1 _13788_ (.A0(_07350_),
    .A1(_07347_),
    .S(net328),
    .X(_07701_));
 sg13g2_o21ai_1 _13789_ (.B1(net53),
    .Y(_07702_),
    .A1(net982),
    .A2(net862));
 sg13g2_a21oi_1 _13790_ (.A1(net804),
    .A2(_07702_),
    .Y(_07703_),
    .B1(net556));
 sg13g2_o21ai_1 _13791_ (.B1(net853),
    .Y(_07704_),
    .A1(net558),
    .A2(_07703_));
 sg13g2_nor3_1 _13792_ (.A(net355),
    .B(_06699_),
    .C(_07704_),
    .Y(_07705_));
 sg13g2_or3_1 _13793_ (.A(_06699_),
    .B(_06685_),
    .C(_07704_),
    .X(_07706_));
 sg13g2_o21ai_1 _13794_ (.B1(_07706_),
    .Y(_07707_),
    .A1(net863),
    .A2(_07704_));
 sg13g2_a221oi_1 _13795_ (.B2(_06687_),
    .C1(_07707_),
    .B1(_07705_),
    .A1(net858),
    .Y(_07708_),
    .A2(_07701_));
 sg13g2_buf_2 fanout325 (.A(net326),
    .X(net325));
 sg13g2_buf_1 fanout324 (.A(_07446_),
    .X(net324));
 sg13g2_nand2_1 _13798_ (.Y(_07711_),
    .A(\dp.rf.rf[19][28] ),
    .B(net807));
 sg13g2_o21ai_1 _13799_ (.B1(_07711_),
    .Y(_01082_),
    .A1(net807),
    .A2(net308));
 sg13g2_o21ai_1 _13800_ (.B1(net54),
    .Y(_07712_),
    .A1(net982),
    .A2(net862));
 sg13g2_a21oi_1 _13801_ (.A1(net804),
    .A2(_07712_),
    .Y(_07713_),
    .B1(net556));
 sg13g2_o21ai_1 _13802_ (.B1(net853),
    .Y(_07714_),
    .A1(net558),
    .A2(_07713_));
 sg13g2_nor4_1 _13803_ (.A(net355),
    .B(_06711_),
    .C(_06721_),
    .D(_07714_),
    .Y(_07715_));
 sg13g2_a22oi_1 _13804_ (.Y(_07716_),
    .B1(_07714_),
    .B2(_06711_),
    .A2(_06725_),
    .A1(net862));
 sg13g2_nor2_1 _13805_ (.A(net328),
    .B(_07360_),
    .Y(_07717_));
 sg13g2_a22oi_1 _13806_ (.Y(_07718_),
    .B1(_07717_),
    .B2(net853),
    .A2(_07358_),
    .A1(net328));
 sg13g2_nor3_1 _13807_ (.A(_07715_),
    .B(_07716_),
    .C(_07718_),
    .Y(_07719_));
 sg13g2_buf_2 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_2 fanout322 (.A(net324),
    .X(net322));
 sg13g2_nand2_1 _13810_ (.Y(_07722_),
    .A(\dp.rf.rf[19][29] ),
    .B(net809));
 sg13g2_o21ai_1 _13811_ (.B1(_07722_),
    .Y(_01083_),
    .A1(net809),
    .A2(net176));
 sg13g2_and2_1 _13812_ (.A(_03826_),
    .B(_07376_),
    .X(_07723_));
 sg13g2_and2_1 _13813_ (.A(_06777_),
    .B(_07373_),
    .X(_07724_));
 sg13g2_o21ai_1 _13814_ (.B1(net56),
    .Y(_07725_),
    .A1(net982),
    .A2(net864));
 sg13g2_a21oi_1 _13815_ (.A1(net804),
    .A2(_07725_),
    .Y(_07726_),
    .B1(net556));
 sg13g2_o21ai_1 _13816_ (.B1(net854),
    .Y(_07727_),
    .A1(net559),
    .A2(_07726_));
 sg13g2_nor4_1 _13817_ (.A(net355),
    .B(_06740_),
    .C(_06744_),
    .D(_07727_),
    .Y(_07728_));
 sg13g2_o21ai_1 _13818_ (.B1(net864),
    .Y(_07729_),
    .A1(_06740_),
    .A2(_06748_));
 sg13g2_nor2b_1 _13819_ (.A(_07727_),
    .B_N(_07729_),
    .Y(_07730_));
 sg13g2_nor4_2 _13820_ (.A(_07723_),
    .B(_07724_),
    .C(_07728_),
    .Y(_07731_),
    .D(_07730_));
 sg13g2_buf_2 fanout321 (.A(net322),
    .X(net321));
 sg13g2_buf_2 fanout320 (.A(net321),
    .X(net320));
 sg13g2_nand2_1 _13823_ (.Y(_07734_),
    .A(\dp.rf.rf[19][30] ),
    .B(net809));
 sg13g2_o21ai_1 _13824_ (.B1(_07734_),
    .Y(_01084_),
    .A1(net809),
    .A2(net173));
 sg13g2_a21oi_1 _13825_ (.A1(_06764_),
    .A2(_06766_),
    .Y(_07735_),
    .B1(net829));
 sg13g2_o21ai_1 _13826_ (.B1(net57),
    .Y(_07736_),
    .A1(net983),
    .A2(net864));
 sg13g2_a21oi_1 _13827_ (.A1(net805),
    .A2(_07736_),
    .Y(_07737_),
    .B1(net557));
 sg13g2_o21ai_1 _13828_ (.B1(net853),
    .Y(_07738_),
    .A1(net559),
    .A2(_07737_));
 sg13g2_a22oi_1 _13829_ (.Y(_07739_),
    .B1(_07738_),
    .B2(_06776_),
    .A2(_07735_),
    .A1(_06763_));
 sg13g2_nor3_1 _13830_ (.A(net1250),
    .B(net933),
    .C(_07385_),
    .Y(_07740_));
 sg13g2_a22oi_1 _13831_ (.Y(_07741_),
    .B1(_07739_),
    .B2(_07740_),
    .A2(_07387_),
    .A1(_03826_));
 sg13g2_buf_2 fanout319 (.A(_07454_),
    .X(net319));
 sg13g2_buf_2 fanout318 (.A(_07454_),
    .X(net318));
 sg13g2_nand2_1 _13834_ (.Y(_07744_),
    .A(\dp.rf.rf[19][31] ),
    .B(net563));
 sg13g2_o21ai_1 _13835_ (.B1(_07744_),
    .Y(_01085_),
    .A1(net563),
    .A2(net167));
 sg13g2_nor2b_1 _13836_ (.A(net1244),
    .B_N(net1256),
    .Y(_07745_));
 sg13g2_and2_1 _13837_ (.A(_05285_),
    .B(_07745_),
    .X(_07746_));
 sg13g2_buf_1 fanout317 (.A(_07454_),
    .X(net317));
 sg13g2_nand2_1 _13839_ (.Y(_07748_),
    .A(_07396_),
    .B(_07746_));
 sg13g2_buf_1 fanout316 (.A(net317),
    .X(net316));
 sg13g2_buf_2 fanout315 (.A(net317),
    .X(net315));
 sg13g2_buf_1 fanout314 (.A(_07468_),
    .X(net314));
 sg13g2_nand2_1 _13843_ (.Y(_07752_),
    .A(\dp.rf.rf[11][0] ),
    .B(net553));
 sg13g2_o21ai_1 _13844_ (.B1(_07752_),
    .Y(_01086_),
    .A1(net300),
    .A2(net553));
 sg13g2_nand2_1 _13845_ (.Y(_07753_),
    .A(\dp.rf.rf[11][1] ),
    .B(net554));
 sg13g2_o21ai_1 _13846_ (.B1(_07753_),
    .Y(_01087_),
    .A1(net296),
    .A2(net554));
 sg13g2_nand2_1 _13847_ (.Y(_07754_),
    .A(\dp.rf.rf[11][2] ),
    .B(net554));
 sg13g2_o21ai_1 _13848_ (.B1(_07754_),
    .Y(_01088_),
    .A1(net320),
    .A2(net554));
 sg13g2_nand2_1 _13849_ (.Y(_07755_),
    .A(\dp.rf.rf[11][3] ),
    .B(net555));
 sg13g2_o21ai_1 _13850_ (.B1(_07755_),
    .Y(_01089_),
    .A1(net317),
    .A2(net555));
 sg13g2_mux2_1 _13851_ (.A0(net294),
    .A1(\dp.rf.rf[11][4] ),
    .S(net553),
    .X(_01090_));
 sg13g2_nand2_1 _13852_ (.Y(_07756_),
    .A(\dp.rf.rf[11][5] ),
    .B(net551));
 sg13g2_o21ai_1 _13853_ (.B1(_07756_),
    .Y(_01091_),
    .A1(net310),
    .A2(net551));
 sg13g2_nand2_1 _13854_ (.Y(_07757_),
    .A(\dp.rf.rf[11][6] ),
    .B(net552));
 sg13g2_o21ai_1 _13855_ (.B1(_07757_),
    .Y(_01092_),
    .A1(net286),
    .A2(net552));
 sg13g2_nand2_1 _13856_ (.Y(_07758_),
    .A(\dp.rf.rf[11][7] ),
    .B(net551));
 sg13g2_o21ai_1 _13857_ (.B1(_07758_),
    .Y(_01093_),
    .A1(net281),
    .A2(net551));
 sg13g2_nand2_1 _13858_ (.Y(_07759_),
    .A(\dp.rf.rf[11][8] ),
    .B(net552));
 sg13g2_o21ai_1 _13859_ (.B1(_07759_),
    .Y(_01094_),
    .A1(net276),
    .A2(net552));
 sg13g2_buf_2 fanout313 (.A(net314),
    .X(net313));
 sg13g2_nand2_1 _13861_ (.Y(_07761_),
    .A(\dp.rf.rf[11][9] ),
    .B(net553));
 sg13g2_o21ai_1 _13862_ (.B1(_07761_),
    .Y(_01095_),
    .A1(net274),
    .A2(net553));
 sg13g2_nand2_1 _13863_ (.Y(_07762_),
    .A(\dp.rf.rf[11][10] ),
    .B(net552));
 sg13g2_o21ai_1 _13864_ (.B1(_07762_),
    .Y(_01096_),
    .A1(net266),
    .A2(net552));
 sg13g2_buf_2 fanout312 (.A(net313),
    .X(net312));
 sg13g2_nand2_1 _13866_ (.Y(_07764_),
    .A(\dp.rf.rf[11][11] ),
    .B(net554));
 sg13g2_o21ai_1 _13867_ (.B1(_07764_),
    .Y(_01097_),
    .A1(net260),
    .A2(net554));
 sg13g2_nand2_1 _13868_ (.Y(_07765_),
    .A(\dp.rf.rf[11][12] ),
    .B(net554));
 sg13g2_o21ai_1 _13869_ (.B1(_07765_),
    .Y(_01098_),
    .A1(net254),
    .A2(net554));
 sg13g2_mux2_1 _13870_ (.A0(net249),
    .A1(\dp.rf.rf[11][13] ),
    .S(net553),
    .X(_01099_));
 sg13g2_nand2_1 _13871_ (.Y(_07766_),
    .A(\dp.rf.rf[11][14] ),
    .B(net546));
 sg13g2_o21ai_1 _13872_ (.B1(_07766_),
    .Y(_01100_),
    .A1(net248),
    .A2(net547));
 sg13g2_nand2_1 _13873_ (.Y(_07767_),
    .A(\dp.rf.rf[11][15] ),
    .B(net551));
 sg13g2_o21ai_1 _13874_ (.B1(_07767_),
    .Y(_01101_),
    .A1(net243),
    .A2(net551));
 sg13g2_nand2_1 _13875_ (.Y(_07768_),
    .A(\dp.rf.rf[11][16] ),
    .B(net551));
 sg13g2_o21ai_1 _13876_ (.B1(_07768_),
    .Y(_01102_),
    .A1(net236),
    .A2(net551));
 sg13g2_nand2_1 _13877_ (.Y(_07769_),
    .A(\dp.rf.rf[11][17] ),
    .B(net547));
 sg13g2_o21ai_1 _13878_ (.B1(_07769_),
    .Y(_01103_),
    .A1(net229),
    .A2(net547));
 sg13g2_nand2_1 _13879_ (.Y(_07770_),
    .A(\dp.rf.rf[11][18] ),
    .B(net553));
 sg13g2_o21ai_1 _13880_ (.B1(_07770_),
    .Y(_01104_),
    .A1(net227),
    .A2(net553));
 sg13g2_nand2_1 _13881_ (.Y(_07771_),
    .A(\dp.rf.rf[11][19] ),
    .B(net547));
 sg13g2_o21ai_1 _13882_ (.B1(_07771_),
    .Y(_01105_),
    .A1(net219),
    .A2(net546));
 sg13g2_buf_2 fanout311 (.A(net314),
    .X(net311));
 sg13g2_nand2_1 _13884_ (.Y(_07773_),
    .A(\dp.rf.rf[11][20] ),
    .B(net549));
 sg13g2_o21ai_1 _13885_ (.B1(_07773_),
    .Y(_01106_),
    .A1(net214),
    .A2(net549));
 sg13g2_nand2_1 _13886_ (.Y(_07774_),
    .A(\dp.rf.rf[11][21] ),
    .B(net548));
 sg13g2_o21ai_1 _13887_ (.B1(_07774_),
    .Y(_01107_),
    .A1(net209),
    .A2(net548));
 sg13g2_buf_2 fanout310 (.A(net314),
    .X(net310));
 sg13g2_nand2_1 _13889_ (.Y(_07776_),
    .A(\dp.rf.rf[11][22] ),
    .B(net549));
 sg13g2_o21ai_1 _13890_ (.B1(_07776_),
    .Y(_01108_),
    .A1(net205),
    .A2(net550));
 sg13g2_nand2_1 _13891_ (.Y(_07777_),
    .A(\dp.rf.rf[11][23] ),
    .B(net546));
 sg13g2_o21ai_1 _13892_ (.B1(_07777_),
    .Y(_01109_),
    .A1(net203),
    .A2(net546));
 sg13g2_nand2_1 _13893_ (.Y(_07778_),
    .A(\dp.rf.rf[11][24] ),
    .B(net548));
 sg13g2_o21ai_1 _13894_ (.B1(_07778_),
    .Y(_01110_),
    .A1(net196),
    .A2(net548));
 sg13g2_nand2_1 _13895_ (.Y(_07779_),
    .A(\dp.rf.rf[11][25] ),
    .B(net548));
 sg13g2_o21ai_1 _13896_ (.B1(_07779_),
    .Y(_01111_),
    .A1(net192),
    .A2(net548));
 sg13g2_nand2_1 _13897_ (.Y(_07780_),
    .A(\dp.rf.rf[11][26] ),
    .B(net549));
 sg13g2_o21ai_1 _13898_ (.B1(_07780_),
    .Y(_01112_),
    .A1(net186),
    .A2(net549));
 sg13g2_nand2_1 _13899_ (.Y(_07781_),
    .A(\dp.rf.rf[11][27] ),
    .B(net546));
 sg13g2_o21ai_1 _13900_ (.B1(_07781_),
    .Y(_01113_),
    .A1(net181),
    .A2(net546));
 sg13g2_nand2_1 _13901_ (.Y(_07782_),
    .A(\dp.rf.rf[11][28] ),
    .B(net548));
 sg13g2_o21ai_1 _13902_ (.B1(_07782_),
    .Y(_01114_),
    .A1(net307),
    .A2(net548));
 sg13g2_nand2_1 _13903_ (.Y(_07783_),
    .A(\dp.rf.rf[11][29] ),
    .B(net549));
 sg13g2_o21ai_1 _13904_ (.B1(_07783_),
    .Y(_01115_),
    .A1(net178),
    .A2(net550));
 sg13g2_buf_1 fanout309 (.A(_07708_),
    .X(net309));
 sg13g2_nand2_1 _13906_ (.Y(_07785_),
    .A(\dp.rf.rf[11][30] ),
    .B(net549));
 sg13g2_o21ai_1 _13907_ (.B1(_07785_),
    .Y(_01116_),
    .A1(net170),
    .A2(net549));
 sg13g2_nand2_1 _13908_ (.Y(_07786_),
    .A(\dp.rf.rf[11][31] ),
    .B(net546));
 sg13g2_o21ai_1 _13909_ (.B1(_07786_),
    .Y(_01117_),
    .A1(net168),
    .A2(net546));
 sg13g2_nand3_1 _13910_ (.B(net1256),
    .C(net1244),
    .A(net1247),
    .Y(_07787_));
 sg13g2_buf_2 fanout308 (.A(net309),
    .X(net308));
 sg13g2_nor2_1 _13912_ (.A(net31),
    .B(_07393_),
    .Y(_07789_));
 sg13g2_nand2_2 _13913_ (.Y(_07790_),
    .A(net1245),
    .B(_07789_));
 sg13g2_buf_2 fanout307 (.A(net308),
    .X(net307));
 sg13g2_nor2_1 _13915_ (.A(_07787_),
    .B(_07790_),
    .Y(_07792_));
 sg13g2_buf_1 fanout306 (.A(net309),
    .X(net306));
 sg13g2_nor2_1 _13917_ (.A(\dp.rf.rf[29][0] ),
    .B(net544),
    .Y(_07794_));
 sg13g2_a21oi_1 _13918_ (.A1(net302),
    .A2(net544),
    .Y(_01118_),
    .B1(_07794_));
 sg13g2_and2_2 _13919_ (.A(net1245),
    .B(_07789_),
    .X(_07795_));
 sg13g2_buf_2 fanout305 (.A(net309),
    .X(net305));
 sg13g2_nand2b_1 _13921_ (.Y(_07797_),
    .B(_07795_),
    .A_N(_07787_));
 sg13g2_buf_1 fanout304 (.A(_07411_),
    .X(net304));
 sg13g2_buf_1 fanout303 (.A(net304),
    .X(net303));
 sg13g2_buf_2 fanout302 (.A(net304),
    .X(net302));
 sg13g2_nand2_1 _13925_ (.Y(_07801_),
    .A(\dp.rf.rf[29][1] ),
    .B(net541));
 sg13g2_o21ai_1 _13926_ (.B1(_07801_),
    .Y(_01119_),
    .A1(net298),
    .A2(net541));
 sg13g2_nand2_1 _13927_ (.Y(_07802_),
    .A(\dp.rf.rf[29][2] ),
    .B(net542));
 sg13g2_o21ai_1 _13928_ (.B1(_07802_),
    .Y(_01120_),
    .A1(net322),
    .A2(net541));
 sg13g2_nand2_1 _13929_ (.Y(_07803_),
    .A(\dp.rf.rf[29][3] ),
    .B(net541));
 sg13g2_o21ai_1 _13930_ (.B1(_07803_),
    .Y(_01121_),
    .A1(net316),
    .A2(net541));
 sg13g2_buf_2 fanout301 (.A(net304),
    .X(net301));
 sg13g2_mux2_1 _13932_ (.A0(\dp.rf.rf[29][4] ),
    .A1(net292),
    .S(net544),
    .X(_01122_));
 sg13g2_nand2_1 _13933_ (.Y(_07805_),
    .A(\dp.rf.rf[29][5] ),
    .B(net539));
 sg13g2_o21ai_1 _13934_ (.B1(_07805_),
    .Y(_01123_),
    .A1(net312),
    .A2(net539));
 sg13g2_nand2_1 _13935_ (.Y(_07806_),
    .A(\dp.rf.rf[29][6] ),
    .B(net540));
 sg13g2_o21ai_1 _13936_ (.B1(_07806_),
    .Y(_01124_),
    .A1(net287),
    .A2(net540));
 sg13g2_buf_2 fanout300 (.A(net301),
    .X(net300));
 sg13g2_nand2_1 _13938_ (.Y(_07808_),
    .A(\dp.rf.rf[29][7] ),
    .B(net540));
 sg13g2_o21ai_1 _13939_ (.B1(_07808_),
    .Y(_01125_),
    .A1(net284),
    .A2(net540));
 sg13g2_nand2_1 _13940_ (.Y(_07809_),
    .A(\dp.rf.rf[29][8] ),
    .B(net542));
 sg13g2_o21ai_1 _13941_ (.B1(_07809_),
    .Y(_01126_),
    .A1(net278),
    .A2(net542));
 sg13g2_nand2_1 _13942_ (.Y(_07810_),
    .A(\dp.rf.rf[29][9] ),
    .B(net539));
 sg13g2_o21ai_1 _13943_ (.B1(_07810_),
    .Y(_01127_),
    .A1(net273),
    .A2(net539));
 sg13g2_nand2_1 _13944_ (.Y(_07811_),
    .A(\dp.rf.rf[29][10] ),
    .B(net541));
 sg13g2_o21ai_1 _13945_ (.B1(_07811_),
    .Y(_01128_),
    .A1(net268),
    .A2(net541));
 sg13g2_nand2_1 _13946_ (.Y(_07812_),
    .A(\dp.rf.rf[29][11] ),
    .B(net542));
 sg13g2_o21ai_1 _13947_ (.B1(_07812_),
    .Y(_01129_),
    .A1(net262),
    .A2(net541));
 sg13g2_buf_1 fanout299 (.A(_07431_),
    .X(net299));
 sg13g2_nand2_1 _13949_ (.Y(_07814_),
    .A(\dp.rf.rf[29][12] ),
    .B(net540));
 sg13g2_o21ai_1 _13950_ (.B1(_07814_),
    .Y(_01130_),
    .A1(net256),
    .A2(net540));
 sg13g2_buf_2 fanout298 (.A(net299),
    .X(net298));
 sg13g2_mux2_1 _13952_ (.A0(\dp.rf.rf[29][13] ),
    .A1(net252),
    .S(net544),
    .X(_01131_));
 sg13g2_nor2_1 _13953_ (.A(\dp.rf.rf[29][14] ),
    .B(net544),
    .Y(_07816_));
 sg13g2_a21oi_1 _13954_ (.A1(net248),
    .A2(net544),
    .Y(_01132_),
    .B1(_07816_));
 sg13g2_nand2_1 _13955_ (.Y(_07817_),
    .A(\dp.rf.rf[29][15] ),
    .B(net539));
 sg13g2_o21ai_1 _13956_ (.B1(_07817_),
    .Y(_01133_),
    .A1(net241),
    .A2(net539));
 sg13g2_nand2_1 _13957_ (.Y(_07818_),
    .A(\dp.rf.rf[29][16] ),
    .B(net539));
 sg13g2_o21ai_1 _13958_ (.B1(_07818_),
    .Y(_01134_),
    .A1(net234),
    .A2(net539));
 sg13g2_nand2_1 _13959_ (.Y(_07819_),
    .A(\dp.rf.rf[29][17] ),
    .B(net538));
 sg13g2_o21ai_1 _13960_ (.B1(_07819_),
    .Y(_01135_),
    .A1(net231),
    .A2(net538));
 sg13g2_nand2_1 _13961_ (.Y(_07820_),
    .A(\dp.rf.rf[29][18] ),
    .B(net537));
 sg13g2_o21ai_1 _13962_ (.B1(_07820_),
    .Y(_01136_),
    .A1(net224),
    .A2(net537));
 sg13g2_buf_2 fanout297 (.A(net299),
    .X(net297));
 sg13g2_nand2_1 _13964_ (.Y(_07822_),
    .A(\dp.rf.rf[29][19] ),
    .B(net537));
 sg13g2_o21ai_1 _13965_ (.B1(_07822_),
    .Y(_01137_),
    .A1(net221),
    .A2(net537));
 sg13g2_nand2_1 _13966_ (.Y(_07823_),
    .A(\dp.rf.rf[29][20] ),
    .B(net538));
 sg13g2_o21ai_1 _13967_ (.B1(_07823_),
    .Y(_01138_),
    .A1(net216),
    .A2(net538));
 sg13g2_nand2_1 _13968_ (.Y(_07824_),
    .A(\dp.rf.rf[29][21] ),
    .B(net536));
 sg13g2_o21ai_1 _13969_ (.B1(_07824_),
    .Y(_01139_),
    .A1(net211),
    .A2(net536));
 sg13g2_buf_1 fanout296 (.A(_07431_),
    .X(net296));
 sg13g2_nor2_1 _13971_ (.A(\dp.rf.rf[29][22] ),
    .B(net545),
    .Y(_07826_));
 sg13g2_a21oi_1 _13972_ (.A1(net208),
    .A2(net545),
    .Y(_01140_),
    .B1(_07826_));
 sg13g2_nand2_1 _13973_ (.Y(_07827_),
    .A(\dp.rf.rf[29][23] ),
    .B(net535));
 sg13g2_o21ai_1 _13974_ (.B1(_07827_),
    .Y(_01141_),
    .A1(net200),
    .A2(net535));
 sg13g2_nand2_1 _13975_ (.Y(_07828_),
    .A(\dp.rf.rf[29][24] ),
    .B(net538));
 sg13g2_o21ai_1 _13976_ (.B1(_07828_),
    .Y(_01142_),
    .A1(net197),
    .A2(net538));
 sg13g2_nand2_1 _13977_ (.Y(_07829_),
    .A(\dp.rf.rf[29][25] ),
    .B(net535));
 sg13g2_o21ai_1 _13978_ (.B1(_07829_),
    .Y(_01143_),
    .A1(net189),
    .A2(net535));
 sg13g2_nand2_1 _13979_ (.Y(_07830_),
    .A(\dp.rf.rf[29][26] ),
    .B(net535));
 sg13g2_o21ai_1 _13980_ (.B1(_07830_),
    .Y(_01144_),
    .A1(net184),
    .A2(net535));
 sg13g2_nand2_1 _13981_ (.Y(_07831_),
    .A(\dp.rf.rf[29][27] ),
    .B(net535));
 sg13g2_o21ai_1 _13982_ (.B1(_07831_),
    .Y(_01145_),
    .A1(net179),
    .A2(net535));
 sg13g2_nand2_1 _13983_ (.Y(_07832_),
    .A(\dp.rf.rf[29][28] ),
    .B(net536));
 sg13g2_o21ai_1 _13984_ (.B1(_07832_),
    .Y(_01146_),
    .A1(net306),
    .A2(net536));
 sg13g2_buf_2 fanout295 (.A(net296),
    .X(net295));
 sg13g2_nor2_1 _13986_ (.A(\dp.rf.rf[29][29] ),
    .B(net544),
    .Y(_07834_));
 sg13g2_a21oi_1 _13987_ (.A1(net174),
    .A2(net545),
    .Y(_01147_),
    .B1(_07834_));
 sg13g2_nor2_1 _13988_ (.A(\dp.rf.rf[29][30] ),
    .B(net544),
    .Y(_07835_));
 sg13g2_a21oi_1 _13989_ (.A1(net173),
    .A2(net545),
    .Y(_01148_),
    .B1(_07835_));
 sg13g2_nand2_1 _13990_ (.Y(_07836_),
    .A(\dp.rf.rf[29][31] ),
    .B(net537));
 sg13g2_o21ai_1 _13991_ (.B1(_07836_),
    .Y(_01149_),
    .A1(net166),
    .A2(net537));
 sg13g2_buf_2 fanout294 (.A(_07462_),
    .X(net294));
 sg13g2_and3_1 _13993_ (.X(_07838_),
    .A(_05285_),
    .B(net1256),
    .C(net1244));
 sg13g2_buf_1 fanout293 (.A(net294),
    .X(net293));
 sg13g2_nor3_2 _13995_ (.A(net1247),
    .B(net1256),
    .C(net1244),
    .Y(_07840_));
 sg13g2_nor4_2 _13996_ (.A(net31),
    .B(net1245),
    .C(_07393_),
    .Y(_07841_),
    .D(_07840_));
 sg13g2_buf_1 fanout292 (.A(net293),
    .X(net292));
 sg13g2_nand2_1 _13998_ (.Y(_07843_),
    .A(_07838_),
    .B(_07841_));
 sg13g2_buf_1 fanout291 (.A(net293),
    .X(net291));
 sg13g2_buf_2 fanout290 (.A(net293),
    .X(net290));
 sg13g2_buf_1 fanout289 (.A(_07476_),
    .X(net289));
 sg13g2_nand2_1 _14002_ (.Y(_07847_),
    .A(\dp.rf.rf[12][0] ),
    .B(net799));
 sg13g2_o21ai_1 _14003_ (.B1(_07847_),
    .Y(_01150_),
    .A1(net300),
    .A2(net796));
 sg13g2_nand2_1 _14004_ (.Y(_07848_),
    .A(\dp.rf.rf[12][1] ),
    .B(net800));
 sg13g2_o21ai_1 _14005_ (.B1(_07848_),
    .Y(_01151_),
    .A1(net295),
    .A2(net800));
 sg13g2_nand2_1 _14006_ (.Y(_07849_),
    .A(\dp.rf.rf[12][2] ),
    .B(net801));
 sg13g2_o21ai_1 _14007_ (.B1(_07849_),
    .Y(_01152_),
    .A1(net320),
    .A2(net801));
 sg13g2_nand2_1 _14008_ (.Y(_07850_),
    .A(\dp.rf.rf[12][3] ),
    .B(net801));
 sg13g2_o21ai_1 _14009_ (.B1(_07850_),
    .Y(_01153_),
    .A1(net315),
    .A2(net801));
 sg13g2_mux2_1 _14010_ (.A0(net291),
    .A1(\dp.rf.rf[12][4] ),
    .S(net796),
    .X(_01154_));
 sg13g2_nand2_1 _14011_ (.Y(_07851_),
    .A(\dp.rf.rf[12][5] ),
    .B(net798));
 sg13g2_o21ai_1 _14012_ (.B1(_07851_),
    .Y(_01155_),
    .A1(net310),
    .A2(net797));
 sg13g2_nand2_1 _14013_ (.Y(_07852_),
    .A(\dp.rf.rf[12][6] ),
    .B(net797));
 sg13g2_o21ai_1 _14014_ (.B1(_07852_),
    .Y(_01156_),
    .A1(net285),
    .A2(net797));
 sg13g2_nand2_1 _14015_ (.Y(_07853_),
    .A(\dp.rf.rf[12][7] ),
    .B(net797));
 sg13g2_o21ai_1 _14016_ (.B1(_07853_),
    .Y(_01157_),
    .A1(net282),
    .A2(net797));
 sg13g2_nand2_1 _14017_ (.Y(_07854_),
    .A(\dp.rf.rf[12][8] ),
    .B(net800));
 sg13g2_o21ai_1 _14018_ (.B1(_07854_),
    .Y(_01158_),
    .A1(net277),
    .A2(net800));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_nand2_1 _14020_ (.Y(_07856_),
    .A(\dp.rf.rf[12][9] ),
    .B(net796));
 sg13g2_o21ai_1 _14021_ (.B1(_07856_),
    .Y(_01159_),
    .A1(net272),
    .A2(net796));
 sg13g2_nand2_1 _14022_ (.Y(_07857_),
    .A(\dp.rf.rf[12][10] ),
    .B(net798));
 sg13g2_o21ai_1 _14023_ (.B1(_07857_),
    .Y(_01160_),
    .A1(net267),
    .A2(net797));
 sg13g2_buf_2 fanout287 (.A(net288),
    .X(net287));
 sg13g2_nand2_1 _14025_ (.Y(_07859_),
    .A(\dp.rf.rf[12][11] ),
    .B(net800));
 sg13g2_o21ai_1 _14026_ (.B1(_07859_),
    .Y(_01161_),
    .A1(net261),
    .A2(net800));
 sg13g2_nand2_1 _14027_ (.Y(_07860_),
    .A(\dp.rf.rf[12][12] ),
    .B(net800));
 sg13g2_o21ai_1 _14028_ (.B1(_07860_),
    .Y(_01162_),
    .A1(net255),
    .A2(net800));
 sg13g2_mux2_1 _14029_ (.A0(net250),
    .A1(\dp.rf.rf[12][13] ),
    .S(net802),
    .X(_01163_));
 sg13g2_buf_2 fanout286 (.A(net289),
    .X(net286));
 sg13g2_nand2_1 _14031_ (.Y(_07862_),
    .A(\dp.rf.rf[12][14] ),
    .B(net793));
 sg13g2_o21ai_1 _14032_ (.B1(_07862_),
    .Y(_01164_),
    .A1(net245),
    .A2(net793));
 sg13g2_nand2_1 _14033_ (.Y(_07863_),
    .A(\dp.rf.rf[12][15] ),
    .B(net797));
 sg13g2_o21ai_1 _14034_ (.B1(_07863_),
    .Y(_01165_),
    .A1(net241),
    .A2(net797));
 sg13g2_nand2_1 _14035_ (.Y(_07864_),
    .A(\dp.rf.rf[12][16] ),
    .B(net798));
 sg13g2_o21ai_1 _14036_ (.B1(_07864_),
    .Y(_01166_),
    .A1(net236),
    .A2(net798));
 sg13g2_nand2_1 _14037_ (.Y(_07865_),
    .A(\dp.rf.rf[12][17] ),
    .B(net795));
 sg13g2_o21ai_1 _14038_ (.B1(_07865_),
    .Y(_01167_),
    .A1(net230),
    .A2(net795));
 sg13g2_nand2_1 _14039_ (.Y(_07866_),
    .A(\dp.rf.rf[12][18] ),
    .B(net796));
 sg13g2_o21ai_1 _14040_ (.B1(_07866_),
    .Y(_01168_),
    .A1(net224),
    .A2(net796));
 sg13g2_nand2_1 _14041_ (.Y(_07867_),
    .A(\dp.rf.rf[12][19] ),
    .B(net796));
 sg13g2_o21ai_1 _14042_ (.B1(_07867_),
    .Y(_01169_),
    .A1(net219),
    .A2(net796));
 sg13g2_buf_2 fanout285 (.A(net289),
    .X(net285));
 sg13g2_nand2_1 _14044_ (.Y(_07869_),
    .A(\dp.rf.rf[12][20] ),
    .B(net794));
 sg13g2_o21ai_1 _14045_ (.B1(_07869_),
    .Y(_01170_),
    .A1(net218),
    .A2(net794));
 sg13g2_nand2_1 _14046_ (.Y(_07870_),
    .A(\dp.rf.rf[12][21] ),
    .B(net792));
 sg13g2_o21ai_1 _14047_ (.B1(_07870_),
    .Y(_01171_),
    .A1(net209),
    .A2(net792));
 sg13g2_buf_2 fanout284 (.A(_07484_),
    .X(net284));
 sg13g2_nand2_1 _14049_ (.Y(_07872_),
    .A(\dp.rf.rf[12][22] ),
    .B(net794));
 sg13g2_o21ai_1 _14050_ (.B1(_07872_),
    .Y(_01172_),
    .A1(net205),
    .A2(net795));
 sg13g2_nand2_1 _14051_ (.Y(_07873_),
    .A(\dp.rf.rf[12][23] ),
    .B(net793));
 sg13g2_o21ai_1 _14052_ (.B1(_07873_),
    .Y(_01173_),
    .A1(net204),
    .A2(net793));
 sg13g2_nand2_1 _14053_ (.Y(_07874_),
    .A(\dp.rf.rf[12][24] ),
    .B(net792));
 sg13g2_o21ai_1 _14054_ (.B1(_07874_),
    .Y(_01174_),
    .A1(net195),
    .A2(net792));
 sg13g2_nand2_1 _14055_ (.Y(_07875_),
    .A(\dp.rf.rf[12][25] ),
    .B(net792));
 sg13g2_o21ai_1 _14056_ (.B1(_07875_),
    .Y(_01175_),
    .A1(net191),
    .A2(net792));
 sg13g2_nand2_1 _14057_ (.Y(_07876_),
    .A(\dp.rf.rf[12][26] ),
    .B(net794));
 sg13g2_o21ai_1 _14058_ (.B1(_07876_),
    .Y(_01176_),
    .A1(net186),
    .A2(net794));
 sg13g2_nand2_1 _14059_ (.Y(_07877_),
    .A(\dp.rf.rf[12][27] ),
    .B(net793));
 sg13g2_o21ai_1 _14060_ (.B1(_07877_),
    .Y(_01177_),
    .A1(net182),
    .A2(net793));
 sg13g2_nand2_1 _14061_ (.Y(_07878_),
    .A(\dp.rf.rf[12][28] ),
    .B(net792));
 sg13g2_o21ai_1 _14062_ (.B1(_07878_),
    .Y(_01178_),
    .A1(net305),
    .A2(net792));
 sg13g2_nand2_1 _14063_ (.Y(_07879_),
    .A(\dp.rf.rf[12][29] ),
    .B(net794));
 sg13g2_o21ai_1 _14064_ (.B1(_07879_),
    .Y(_01179_),
    .A1(net177),
    .A2(net795));
 sg13g2_nand2_1 _14065_ (.Y(_07880_),
    .A(\dp.rf.rf[12][30] ),
    .B(net794));
 sg13g2_o21ai_1 _14066_ (.B1(_07880_),
    .Y(_01180_),
    .A1(net171),
    .A2(net794));
 sg13g2_nand2_1 _14067_ (.Y(_07881_),
    .A(\dp.rf.rf[12][31] ),
    .B(net793));
 sg13g2_o21ai_1 _14068_ (.B1(_07881_),
    .Y(_01181_),
    .A1(net167),
    .A2(net793));
 sg13g2_nand2_1 _14069_ (.Y(_07882_),
    .A(_07795_),
    .B(_07838_));
 sg13g2_buf_2 fanout283 (.A(net284),
    .X(net283));
 sg13g2_buf_2 fanout282 (.A(_07484_),
    .X(net282));
 sg13g2_buf_2 fanout281 (.A(net282),
    .X(net281));
 sg13g2_nand2_1 _14073_ (.Y(_07886_),
    .A(\dp.rf.rf[13][0] ),
    .B(net531));
 sg13g2_o21ai_1 _14074_ (.B1(_07886_),
    .Y(_01182_),
    .A1(net301),
    .A2(net531));
 sg13g2_nand2_1 _14075_ (.Y(_07887_),
    .A(\dp.rf.rf[13][1] ),
    .B(net532));
 sg13g2_o21ai_1 _14076_ (.B1(_07887_),
    .Y(_01183_),
    .A1(net295),
    .A2(net532));
 sg13g2_nand2_1 _14077_ (.Y(_07888_),
    .A(\dp.rf.rf[13][2] ),
    .B(net533));
 sg13g2_o21ai_1 _14078_ (.B1(_07888_),
    .Y(_01184_),
    .A1(net321),
    .A2(net532));
 sg13g2_buf_1 fanout280 (.A(_07498_),
    .X(net280));
 sg13g2_nand2_1 _14080_ (.Y(_07890_),
    .A(\dp.rf.rf[13][3] ),
    .B(net533));
 sg13g2_o21ai_1 _14081_ (.B1(_07890_),
    .Y(_01185_),
    .A1(net317),
    .A2(net532));
 sg13g2_nand3_1 _14082_ (.B(net1256),
    .C(net1244),
    .A(_05285_),
    .Y(_07891_));
 sg13g2_nor2_2 _14083_ (.A(_07790_),
    .B(_07891_),
    .Y(_07892_));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_mux2_1 _14085_ (.A0(\dp.rf.rf[13][4] ),
    .A1(net290),
    .S(_07892_),
    .X(_01186_));
 sg13g2_nand2_1 _14086_ (.Y(_07894_),
    .A(\dp.rf.rf[13][5] ),
    .B(net529));
 sg13g2_o21ai_1 _14087_ (.B1(_07894_),
    .Y(_01187_),
    .A1(net310),
    .A2(net529));
 sg13g2_nand2_1 _14088_ (.Y(_07895_),
    .A(\dp.rf.rf[13][6] ),
    .B(net529));
 sg13g2_o21ai_1 _14089_ (.B1(_07895_),
    .Y(_01188_),
    .A1(net285),
    .A2(net529));
 sg13g2_nand2_1 _14090_ (.Y(_07896_),
    .A(\dp.rf.rf[13][7] ),
    .B(net530));
 sg13g2_o21ai_1 _14091_ (.B1(_07896_),
    .Y(_01189_),
    .A1(net282),
    .A2(net530));
 sg13g2_nand2_1 _14092_ (.Y(_07897_),
    .A(\dp.rf.rf[13][8] ),
    .B(net530));
 sg13g2_o21ai_1 _14093_ (.B1(_07897_),
    .Y(_01190_),
    .A1(net276),
    .A2(net530));
 sg13g2_nand2_1 _14094_ (.Y(_07898_),
    .A(\dp.rf.rf[13][9] ),
    .B(net531));
 sg13g2_o21ai_1 _14095_ (.B1(_07898_),
    .Y(_01191_),
    .A1(net272),
    .A2(net531));
 sg13g2_nand2_1 _14096_ (.Y(_07899_),
    .A(\dp.rf.rf[13][10] ),
    .B(net530));
 sg13g2_o21ai_1 _14097_ (.B1(_07899_),
    .Y(_01192_),
    .A1(net266),
    .A2(net530));
 sg13g2_buf_2 fanout278 (.A(net279),
    .X(net278));
 sg13g2_nand2_1 _14099_ (.Y(_07901_),
    .A(\dp.rf.rf[13][11] ),
    .B(net532));
 sg13g2_o21ai_1 _14100_ (.B1(_07901_),
    .Y(_01193_),
    .A1(net260),
    .A2(net532));
 sg13g2_nand2_1 _14101_ (.Y(_07902_),
    .A(\dp.rf.rf[13][12] ),
    .B(net532));
 sg13g2_o21ai_1 _14102_ (.B1(_07902_),
    .Y(_01194_),
    .A1(net254),
    .A2(net532));
 sg13g2_mux2_1 _14103_ (.A0(\dp.rf.rf[13][13] ),
    .A1(net249),
    .S(_07892_),
    .X(_01195_));
 sg13g2_nor2_1 _14104_ (.A(\dp.rf.rf[13][14] ),
    .B(_07892_),
    .Y(_07903_));
 sg13g2_a21oi_1 _14105_ (.A1(net246),
    .A2(_07892_),
    .Y(_01196_),
    .B1(_07903_));
 sg13g2_nand2_1 _14106_ (.Y(_07904_),
    .A(\dp.rf.rf[13][15] ),
    .B(net529));
 sg13g2_o21ai_1 _14107_ (.B1(_07904_),
    .Y(_01197_),
    .A1(net242),
    .A2(net529));
 sg13g2_buf_2 fanout277 (.A(net280),
    .X(net277));
 sg13g2_nand2_1 _14109_ (.Y(_07906_),
    .A(\dp.rf.rf[13][16] ),
    .B(net529));
 sg13g2_o21ai_1 _14110_ (.B1(_07906_),
    .Y(_01198_),
    .A1(net236),
    .A2(net529));
 sg13g2_buf_2 fanout276 (.A(net280),
    .X(net276));
 sg13g2_nand2_1 _14112_ (.Y(_07908_),
    .A(\dp.rf.rf[13][17] ),
    .B(net528));
 sg13g2_o21ai_1 _14113_ (.B1(_07908_),
    .Y(_01199_),
    .A1(net230),
    .A2(net528));
 sg13g2_nand2_1 _14114_ (.Y(_07909_),
    .A(\dp.rf.rf[13][18] ),
    .B(net531));
 sg13g2_o21ai_1 _14115_ (.B1(_07909_),
    .Y(_01200_),
    .A1(net226),
    .A2(net531));
 sg13g2_nand2_1 _14116_ (.Y(_07910_),
    .A(\dp.rf.rf[13][19] ),
    .B(net531));
 sg13g2_o21ai_1 _14117_ (.B1(_07910_),
    .Y(_01201_),
    .A1(net219),
    .A2(net531));
 sg13g2_buf_1 fanout275 (.A(_07507_),
    .X(net275));
 sg13g2_nand2_1 _14119_ (.Y(_07912_),
    .A(\dp.rf.rf[13][20] ),
    .B(net528));
 sg13g2_o21ai_1 _14120_ (.B1(_07912_),
    .Y(_01202_),
    .A1(net215),
    .A2(net528));
 sg13g2_nand2_1 _14121_ (.Y(_07913_),
    .A(\dp.rf.rf[13][21] ),
    .B(net526));
 sg13g2_o21ai_1 _14122_ (.B1(_07913_),
    .Y(_01203_),
    .A1(net210),
    .A2(net526));
 sg13g2_nor2_1 _14123_ (.A(\dp.rf.rf[13][22] ),
    .B(_07892_),
    .Y(_07914_));
 sg13g2_a21oi_1 _14124_ (.A1(net205),
    .A2(_07892_),
    .Y(_01204_),
    .B1(_07914_));
 sg13g2_nand2_1 _14125_ (.Y(_07915_),
    .A(\dp.rf.rf[13][23] ),
    .B(net527));
 sg13g2_o21ai_1 _14126_ (.B1(_07915_),
    .Y(_01205_),
    .A1(net203),
    .A2(net527));
 sg13g2_nand2_1 _14127_ (.Y(_07916_),
    .A(\dp.rf.rf[13][24] ),
    .B(net526));
 sg13g2_o21ai_1 _14128_ (.B1(_07916_),
    .Y(_01206_),
    .A1(net195),
    .A2(net526));
 sg13g2_nand2_1 _14129_ (.Y(_07917_),
    .A(\dp.rf.rf[13][25] ),
    .B(net526));
 sg13g2_o21ai_1 _14130_ (.B1(_07917_),
    .Y(_01207_),
    .A1(net191),
    .A2(net526));
 sg13g2_nand2_1 _14131_ (.Y(_07918_),
    .A(\dp.rf.rf[13][26] ),
    .B(net534));
 sg13g2_o21ai_1 _14132_ (.B1(_07918_),
    .Y(_01208_),
    .A1(net187),
    .A2(net534));
 sg13g2_nand2_1 _14133_ (.Y(_07919_),
    .A(\dp.rf.rf[13][27] ),
    .B(net527));
 sg13g2_o21ai_1 _14134_ (.B1(_07919_),
    .Y(_01209_),
    .A1(net181),
    .A2(net527));
 sg13g2_nand2_1 _14135_ (.Y(_07920_),
    .A(\dp.rf.rf[13][28] ),
    .B(net526));
 sg13g2_o21ai_1 _14136_ (.B1(_07920_),
    .Y(_01210_),
    .A1(net305),
    .A2(net526));
 sg13g2_nor2_1 _14137_ (.A(\dp.rf.rf[13][29] ),
    .B(_07892_),
    .Y(_07921_));
 sg13g2_a21oi_1 _14138_ (.A1(net177),
    .A2(_07892_),
    .Y(_01211_),
    .B1(_07921_));
 sg13g2_nand2_1 _14139_ (.Y(_07922_),
    .A(\dp.rf.rf[13][30] ),
    .B(net528));
 sg13g2_o21ai_1 _14140_ (.B1(_07922_),
    .Y(_01212_),
    .A1(net170),
    .A2(net528));
 sg13g2_nand2_1 _14141_ (.Y(_07923_),
    .A(\dp.rf.rf[13][31] ),
    .B(net527));
 sg13g2_o21ai_1 _14142_ (.B1(_07923_),
    .Y(_01213_),
    .A1(net167),
    .A2(net527));
 sg13g2_nand2b_2 _14143_ (.Y(_07924_),
    .B(_07395_),
    .A_N(net1246));
 sg13g2_buf_2 fanout274 (.A(_07507_),
    .X(net274));
 sg13g2_nor2_1 _14145_ (.A(_07891_),
    .B(_07924_),
    .Y(_07926_));
 sg13g2_buf_1 fanout273 (.A(_07507_),
    .X(net273));
 sg13g2_buf_2 fanout272 (.A(net273),
    .X(net272));
 sg13g2_nor2_1 _14148_ (.A(\dp.rf.rf[14][0] ),
    .B(net525),
    .Y(_07929_));
 sg13g2_a21oi_1 _14149_ (.A1(net304),
    .A2(net525),
    .Y(_01214_),
    .B1(_07929_));
 sg13g2_nor3_2 _14150_ (.A(_05645_),
    .B(net1246),
    .C(_07393_),
    .Y(_07930_));
 sg13g2_buf_2 fanout271 (.A(net273),
    .X(net271));
 sg13g2_nand2_1 _14152_ (.Y(_07932_),
    .A(_07838_),
    .B(_07930_));
 sg13g2_buf_1 fanout270 (.A(_07516_),
    .X(net270));
 sg13g2_buf_2 fanout269 (.A(net270),
    .X(net269));
 sg13g2_buf_2 fanout268 (.A(net269),
    .X(net268));
 sg13g2_buf_1 fanout267 (.A(net270),
    .X(net267));
 sg13g2_nand2_1 _14157_ (.Y(_07937_),
    .A(\dp.rf.rf[14][1] ),
    .B(net789));
 sg13g2_o21ai_1 _14158_ (.B1(_07937_),
    .Y(_01215_),
    .A1(net295),
    .A2(net789));
 sg13g2_nand2_1 _14159_ (.Y(_07938_),
    .A(\dp.rf.rf[14][2] ),
    .B(net790));
 sg13g2_o21ai_1 _14160_ (.B1(_07938_),
    .Y(_01216_),
    .A1(net320),
    .A2(net789));
 sg13g2_nand2_1 _14161_ (.Y(_07939_),
    .A(\dp.rf.rf[14][3] ),
    .B(net790));
 sg13g2_o21ai_1 _14162_ (.B1(_07939_),
    .Y(_01217_),
    .A1(net315),
    .A2(net790));
 sg13g2_mux2_1 _14163_ (.A0(\dp.rf.rf[14][4] ),
    .A1(net291),
    .S(net525),
    .X(_01218_));
 sg13g2_nand2_1 _14164_ (.Y(_07940_),
    .A(\dp.rf.rf[14][5] ),
    .B(net786));
 sg13g2_o21ai_1 _14165_ (.B1(_07940_),
    .Y(_01219_),
    .A1(net310),
    .A2(net786));
 sg13g2_nand2_1 _14166_ (.Y(_07941_),
    .A(\dp.rf.rf[14][6] ),
    .B(net786));
 sg13g2_o21ai_1 _14167_ (.B1(_07941_),
    .Y(_01220_),
    .A1(net285),
    .A2(net786));
 sg13g2_nand2_1 _14168_ (.Y(_07942_),
    .A(\dp.rf.rf[14][7] ),
    .B(net787));
 sg13g2_o21ai_1 _14169_ (.B1(_07942_),
    .Y(_01221_),
    .A1(net282),
    .A2(net786));
 sg13g2_buf_2 fanout266 (.A(net270),
    .X(net266));
 sg13g2_nand2_1 _14171_ (.Y(_07944_),
    .A(\dp.rf.rf[14][8] ),
    .B(net789));
 sg13g2_o21ai_1 _14172_ (.B1(_07944_),
    .Y(_01222_),
    .A1(net277),
    .A2(net789));
 sg13g2_nand2_1 _14173_ (.Y(_07945_),
    .A(\dp.rf.rf[14][9] ),
    .B(net788));
 sg13g2_o21ai_1 _14174_ (.B1(_07945_),
    .Y(_01223_),
    .A1(net272),
    .A2(net788));
 sg13g2_nand2_1 _14175_ (.Y(_07946_),
    .A(\dp.rf.rf[14][10] ),
    .B(net787));
 sg13g2_o21ai_1 _14176_ (.B1(_07946_),
    .Y(_01224_),
    .A1(net267),
    .A2(net787));
 sg13g2_nand2_1 _14177_ (.Y(_07947_),
    .A(\dp.rf.rf[14][11] ),
    .B(net790));
 sg13g2_o21ai_1 _14178_ (.B1(_07947_),
    .Y(_01225_),
    .A1(net261),
    .A2(net789));
 sg13g2_buf_1 fanout265 (.A(_07526_),
    .X(net265));
 sg13g2_nand2_1 _14180_ (.Y(_07949_),
    .A(\dp.rf.rf[14][12] ),
    .B(net789));
 sg13g2_o21ai_1 _14181_ (.B1(_07949_),
    .Y(_01226_),
    .A1(net255),
    .A2(net789));
 sg13g2_mux2_1 _14182_ (.A0(\dp.rf.rf[14][13] ),
    .A1(net249),
    .S(net525),
    .X(_01227_));
 sg13g2_nor2_1 _14183_ (.A(\dp.rf.rf[14][14] ),
    .B(net524),
    .Y(_07950_));
 sg13g2_a21oi_1 _14184_ (.A1(_07550_),
    .A2(net524),
    .Y(_01228_),
    .B1(_07950_));
 sg13g2_nand2_1 _14185_ (.Y(_07951_),
    .A(\dp.rf.rf[14][15] ),
    .B(net786));
 sg13g2_o21ai_1 _14186_ (.B1(_07951_),
    .Y(_01229_),
    .A1(net241),
    .A2(net786));
 sg13g2_nand2_1 _14187_ (.Y(_07952_),
    .A(\dp.rf.rf[14][16] ),
    .B(net787));
 sg13g2_o21ai_1 _14188_ (.B1(_07952_),
    .Y(_01230_),
    .A1(net236),
    .A2(net786));
 sg13g2_nand2_1 _14189_ (.Y(_07953_),
    .A(\dp.rf.rf[14][17] ),
    .B(net785));
 sg13g2_o21ai_1 _14190_ (.B1(_07953_),
    .Y(_01231_),
    .A1(net230),
    .A2(net785));
 sg13g2_nand2_1 _14191_ (.Y(_07954_),
    .A(\dp.rf.rf[14][18] ),
    .B(net788));
 sg13g2_o21ai_1 _14192_ (.B1(_07954_),
    .Y(_01232_),
    .A1(net225),
    .A2(net788));
 sg13g2_nand2_1 _14193_ (.Y(_07955_),
    .A(\dp.rf.rf[14][19] ),
    .B(net788));
 sg13g2_o21ai_1 _14194_ (.B1(_07955_),
    .Y(_01233_),
    .A1(net219),
    .A2(net788));
 sg13g2_nor2_1 _14195_ (.A(\dp.rf.rf[14][20] ),
    .B(net524),
    .Y(_07956_));
 sg13g2_a21oi_1 _14196_ (.A1(net215),
    .A2(net524),
    .Y(_01234_),
    .B1(_07956_));
 sg13g2_nand2_1 _14197_ (.Y(_07957_),
    .A(\dp.rf.rf[14][21] ),
    .B(net783));
 sg13g2_o21ai_1 _14198_ (.B1(_07957_),
    .Y(_01235_),
    .A1(net209),
    .A2(net784));
 sg13g2_nor2_1 _14199_ (.A(\dp.rf.rf[14][22] ),
    .B(net524),
    .Y(_07958_));
 sg13g2_a21oi_1 _14200_ (.A1(net206),
    .A2(net525),
    .Y(_01236_),
    .B1(_07958_));
 sg13g2_nand2_1 _14201_ (.Y(_07959_),
    .A(\dp.rf.rf[14][23] ),
    .B(net784));
 sg13g2_o21ai_1 _14202_ (.B1(_07959_),
    .Y(_01237_),
    .A1(net204),
    .A2(net784));
 sg13g2_nand2_1 _14203_ (.Y(_07960_),
    .A(\dp.rf.rf[14][24] ),
    .B(net783));
 sg13g2_o21ai_1 _14204_ (.B1(_07960_),
    .Y(_01238_),
    .A1(net195),
    .A2(net784));
 sg13g2_nand2_1 _14205_ (.Y(_07961_),
    .A(\dp.rf.rf[14][25] ),
    .B(net783));
 sg13g2_o21ai_1 _14206_ (.B1(_07961_),
    .Y(_01239_),
    .A1(net191),
    .A2(net783));
 sg13g2_nand2_1 _14207_ (.Y(_07962_),
    .A(\dp.rf.rf[14][26] ),
    .B(net785));
 sg13g2_o21ai_1 _14208_ (.B1(_07962_),
    .Y(_01240_),
    .A1(net186),
    .A2(net785));
 sg13g2_nand2_1 _14209_ (.Y(_07963_),
    .A(\dp.rf.rf[14][27] ),
    .B(net783));
 sg13g2_o21ai_1 _14210_ (.B1(_07963_),
    .Y(_01241_),
    .A1(net181),
    .A2(net783));
 sg13g2_nand2_1 _14211_ (.Y(_07964_),
    .A(\dp.rf.rf[14][28] ),
    .B(net783));
 sg13g2_o21ai_1 _14212_ (.B1(_07964_),
    .Y(_01242_),
    .A1(net305),
    .A2(net783));
 sg13g2_nor2_1 _14213_ (.A(\dp.rf.rf[14][29] ),
    .B(net524),
    .Y(_07965_));
 sg13g2_a21oi_1 _14214_ (.A1(net177),
    .A2(net525),
    .Y(_01243_),
    .B1(_07965_));
 sg13g2_nor2_1 _14215_ (.A(\dp.rf.rf[14][30] ),
    .B(net524),
    .Y(_07966_));
 sg13g2_a21oi_1 _14216_ (.A1(net171),
    .A2(net524),
    .Y(_01244_),
    .B1(_07966_));
 sg13g2_nand2_1 _14217_ (.Y(_07967_),
    .A(\dp.rf.rf[14][31] ),
    .B(net784));
 sg13g2_o21ai_1 _14218_ (.B1(_07967_),
    .Y(_01245_),
    .A1(net166),
    .A2(net784));
 sg13g2_nand2_1 _14219_ (.Y(_07968_),
    .A(_07396_),
    .B(_07838_));
 sg13g2_buf_1 fanout264 (.A(net265),
    .X(net264));
 sg13g2_buf_2 fanout263 (.A(net265),
    .X(net263));
 sg13g2_buf_2 fanout262 (.A(net265),
    .X(net262));
 sg13g2_nand2_1 _14223_ (.Y(_07972_),
    .A(\dp.rf.rf[15][0] ),
    .B(net518));
 sg13g2_o21ai_1 _14224_ (.B1(_07972_),
    .Y(_01246_),
    .A1(net300),
    .A2(net518));
 sg13g2_nand2_1 _14225_ (.Y(_07973_),
    .A(\dp.rf.rf[15][1] ),
    .B(net522));
 sg13g2_o21ai_1 _14226_ (.B1(_07973_),
    .Y(_01247_),
    .A1(net295),
    .A2(net522));
 sg13g2_nand2_1 _14227_ (.Y(_07974_),
    .A(\dp.rf.rf[15][2] ),
    .B(net523));
 sg13g2_o21ai_1 _14228_ (.B1(_07974_),
    .Y(_01248_),
    .A1(net321),
    .A2(net523));
 sg13g2_nand2_1 _14229_ (.Y(_07975_),
    .A(\dp.rf.rf[15][3] ),
    .B(net522));
 sg13g2_o21ai_1 _14230_ (.B1(_07975_),
    .Y(_01249_),
    .A1(net317),
    .A2(net522));
 sg13g2_mux2_1 _14231_ (.A0(net291),
    .A1(\dp.rf.rf[15][4] ),
    .S(net521),
    .X(_01250_));
 sg13g2_nand2_1 _14232_ (.Y(_07976_),
    .A(\dp.rf.rf[15][5] ),
    .B(net519));
 sg13g2_o21ai_1 _14233_ (.B1(_07976_),
    .Y(_01251_),
    .A1(net310),
    .A2(net519));
 sg13g2_nand2_1 _14234_ (.Y(_07977_),
    .A(\dp.rf.rf[15][6] ),
    .B(net519));
 sg13g2_o21ai_1 _14235_ (.B1(_07977_),
    .Y(_01252_),
    .A1(net285),
    .A2(net519));
 sg13g2_nand2_1 _14236_ (.Y(_07978_),
    .A(\dp.rf.rf[15][7] ),
    .B(net520));
 sg13g2_o21ai_1 _14237_ (.B1(_07978_),
    .Y(_01253_),
    .A1(net282),
    .A2(net520));
 sg13g2_nand2_1 _14238_ (.Y(_07979_),
    .A(\dp.rf.rf[15][8] ),
    .B(net520));
 sg13g2_o21ai_1 _14239_ (.B1(_07979_),
    .Y(_01254_),
    .A1(net277),
    .A2(net520));
 sg13g2_buf_1 fanout261 (.A(net262),
    .X(net261));
 sg13g2_nand2_1 _14241_ (.Y(_07981_),
    .A(\dp.rf.rf[15][9] ),
    .B(net518));
 sg13g2_o21ai_1 _14242_ (.B1(_07981_),
    .Y(_01255_),
    .A1(net274),
    .A2(net518));
 sg13g2_nand2_1 _14243_ (.Y(_07982_),
    .A(\dp.rf.rf[15][10] ),
    .B(net520));
 sg13g2_o21ai_1 _14244_ (.B1(_07982_),
    .Y(_01256_),
    .A1(net267),
    .A2(net520));
 sg13g2_buf_2 fanout260 (.A(net261),
    .X(net260));
 sg13g2_nand2_1 _14246_ (.Y(_07984_),
    .A(\dp.rf.rf[15][11] ),
    .B(net522));
 sg13g2_o21ai_1 _14247_ (.B1(_07984_),
    .Y(_01257_),
    .A1(net261),
    .A2(net522));
 sg13g2_nand2_1 _14248_ (.Y(_07985_),
    .A(\dp.rf.rf[15][12] ),
    .B(net522));
 sg13g2_o21ai_1 _14249_ (.B1(_07985_),
    .Y(_01258_),
    .A1(net255),
    .A2(net522));
 sg13g2_mux2_1 _14250_ (.A0(net249),
    .A1(\dp.rf.rf[15][13] ),
    .S(net521),
    .X(_01259_));
 sg13g2_nand2_1 _14251_ (.Y(_07986_),
    .A(\dp.rf.rf[15][14] ),
    .B(net515));
 sg13g2_o21ai_1 _14252_ (.B1(_07986_),
    .Y(_01260_),
    .A1(net246),
    .A2(net515));
 sg13g2_nand2_1 _14253_ (.Y(_07987_),
    .A(\dp.rf.rf[15][15] ),
    .B(net519));
 sg13g2_o21ai_1 _14254_ (.B1(_07987_),
    .Y(_01261_),
    .A1(net243),
    .A2(net519));
 sg13g2_nand2_1 _14255_ (.Y(_07988_),
    .A(\dp.rf.rf[15][16] ),
    .B(net519));
 sg13g2_o21ai_1 _14256_ (.B1(_07988_),
    .Y(_01262_),
    .A1(net236),
    .A2(net519));
 sg13g2_nand2_1 _14257_ (.Y(_07989_),
    .A(\dp.rf.rf[15][17] ),
    .B(net515));
 sg13g2_o21ai_1 _14258_ (.B1(_07989_),
    .Y(_01263_),
    .A1(net230),
    .A2(net515));
 sg13g2_nand2_1 _14259_ (.Y(_07990_),
    .A(\dp.rf.rf[15][18] ),
    .B(net518));
 sg13g2_o21ai_1 _14260_ (.B1(_07990_),
    .Y(_01264_),
    .A1(net225),
    .A2(net518));
 sg13g2_nand2_1 _14261_ (.Y(_07991_),
    .A(\dp.rf.rf[15][19] ),
    .B(net518));
 sg13g2_o21ai_1 _14262_ (.B1(_07991_),
    .Y(_01265_),
    .A1(net219),
    .A2(net518));
 sg13g2_buf_1 fanout259 (.A(_07534_),
    .X(net259));
 sg13g2_nand2_1 _14264_ (.Y(_07993_),
    .A(\dp.rf.rf[15][20] ),
    .B(net516));
 sg13g2_o21ai_1 _14265_ (.B1(_07993_),
    .Y(_01266_),
    .A1(net215),
    .A2(net516));
 sg13g2_nand2_1 _14266_ (.Y(_07994_),
    .A(\dp.rf.rf[15][21] ),
    .B(net515));
 sg13g2_o21ai_1 _14267_ (.B1(_07994_),
    .Y(_01267_),
    .A1(net209),
    .A2(net514));
 sg13g2_buf_1 fanout258 (.A(net259),
    .X(net258));
 sg13g2_nand2_1 _14269_ (.Y(_07996_),
    .A(\dp.rf.rf[15][22] ),
    .B(net516));
 sg13g2_o21ai_1 _14270_ (.B1(_07996_),
    .Y(_01268_),
    .A1(net206),
    .A2(net517));
 sg13g2_nand2_1 _14271_ (.Y(_07997_),
    .A(\dp.rf.rf[15][23] ),
    .B(net515));
 sg13g2_o21ai_1 _14272_ (.B1(_07997_),
    .Y(_01269_),
    .A1(net202),
    .A2(net517));
 sg13g2_nand2_1 _14273_ (.Y(_07998_),
    .A(\dp.rf.rf[15][24] ),
    .B(net514));
 sg13g2_o21ai_1 _14274_ (.B1(_07998_),
    .Y(_01270_),
    .A1(net195),
    .A2(net515));
 sg13g2_nand2_1 _14275_ (.Y(_07999_),
    .A(\dp.rf.rf[15][25] ),
    .B(net514));
 sg13g2_o21ai_1 _14276_ (.B1(_07999_),
    .Y(_01271_),
    .A1(net192),
    .A2(net514));
 sg13g2_nand2_1 _14277_ (.Y(_08000_),
    .A(\dp.rf.rf[15][26] ),
    .B(net516));
 sg13g2_o21ai_1 _14278_ (.B1(_08000_),
    .Y(_01272_),
    .A1(net186),
    .A2(net516));
 sg13g2_nand2_1 _14279_ (.Y(_08001_),
    .A(\dp.rf.rf[15][27] ),
    .B(net514));
 sg13g2_o21ai_1 _14280_ (.B1(_08001_),
    .Y(_01273_),
    .A1(net182),
    .A2(net514));
 sg13g2_nand2_1 _14281_ (.Y(_08002_),
    .A(\dp.rf.rf[15][28] ),
    .B(net514));
 sg13g2_o21ai_1 _14282_ (.B1(_08002_),
    .Y(_01274_),
    .A1(net305),
    .A2(net514));
 sg13g2_nand2_1 _14283_ (.Y(_08003_),
    .A(\dp.rf.rf[15][29] ),
    .B(net516));
 sg13g2_o21ai_1 _14284_ (.B1(_08003_),
    .Y(_01275_),
    .A1(net177),
    .A2(net517));
 sg13g2_nand2_1 _14285_ (.Y(_08004_),
    .A(\dp.rf.rf[15][30] ),
    .B(net516));
 sg13g2_o21ai_1 _14286_ (.B1(_08004_),
    .Y(_01276_),
    .A1(net170),
    .A2(net516));
 sg13g2_nand2_1 _14287_ (.Y(_08005_),
    .A(\dp.rf.rf[15][31] ),
    .B(net517));
 sg13g2_o21ai_1 _14288_ (.B1(_08005_),
    .Y(_01277_),
    .A1(net169),
    .A2(net517));
 sg13g2_nand2_1 _14289_ (.Y(_08006_),
    .A(_07390_),
    .B(_07841_));
 sg13g2_buf_1 fanout257 (.A(net258),
    .X(net257));
 sg13g2_buf_2 fanout256 (.A(net258),
    .X(net256));
 sg13g2_buf_1 fanout255 (.A(_07534_),
    .X(net255));
 sg13g2_nand2_1 _14293_ (.Y(_08010_),
    .A(\dp.rf.rf[16][0] ),
    .B(net779));
 sg13g2_o21ai_1 _14294_ (.B1(_08010_),
    .Y(_01278_),
    .A1(net303),
    .A2(net779));
 sg13g2_nand2_1 _14295_ (.Y(_08011_),
    .A(\dp.rf.rf[16][1] ),
    .B(net782));
 sg13g2_o21ai_1 _14296_ (.B1(_08011_),
    .Y(_01279_),
    .A1(net297),
    .A2(net782));
 sg13g2_nand2_1 _14297_ (.Y(_08012_),
    .A(\dp.rf.rf[16][2] ),
    .B(net781));
 sg13g2_o21ai_1 _14298_ (.B1(_08012_),
    .Y(_01280_),
    .A1(net323),
    .A2(net781));
 sg13g2_nand2_1 _14299_ (.Y(_08013_),
    .A(\dp.rf.rf[16][3] ),
    .B(net781));
 sg13g2_o21ai_1 _14300_ (.B1(_08013_),
    .Y(_01281_),
    .A1(net319),
    .A2(net781));
 sg13g2_buf_2 fanout254 (.A(net255),
    .X(net254));
 sg13g2_nand2_1 _14302_ (.Y(_08015_),
    .A(net1247),
    .B(_07389_));
 sg13g2_or4_2 _14303_ (.A(net31),
    .B(net1246),
    .C(_07393_),
    .D(_07840_),
    .X(_08016_));
 sg13g2_buf_1 fanout253 (.A(_07543_),
    .X(net253));
 sg13g2_nor2_1 _14305_ (.A(_08015_),
    .B(_08016_),
    .Y(_08018_));
 sg13g2_buf_2 fanout252 (.A(net253),
    .X(net252));
 sg13g2_mux2_1 _14307_ (.A0(\dp.rf.rf[16][4] ),
    .A1(net290),
    .S(net773),
    .X(_01282_));
 sg13g2_nand2_1 _14308_ (.Y(_08020_),
    .A(\dp.rf.rf[16][5] ),
    .B(net780));
 sg13g2_o21ai_1 _14309_ (.B1(_08020_),
    .Y(_01283_),
    .A1(net312),
    .A2(net780));
 sg13g2_buf_2 fanout251 (.A(net252),
    .X(net251));
 sg13g2_nand2_1 _14311_ (.Y(_08022_),
    .A(\dp.rf.rf[16][6] ),
    .B(net782));
 sg13g2_o21ai_1 _14312_ (.B1(_08022_),
    .Y(_01284_),
    .A1(net288),
    .A2(net782));
 sg13g2_nand2_1 _14313_ (.Y(_08023_),
    .A(\dp.rf.rf[16][7] ),
    .B(net779));
 sg13g2_o21ai_1 _14314_ (.B1(_08023_),
    .Y(_01285_),
    .A1(_07484_),
    .A2(net779));
 sg13g2_nand2_1 _14315_ (.Y(_08024_),
    .A(\dp.rf.rf[16][8] ),
    .B(net781));
 sg13g2_o21ai_1 _14316_ (.B1(_08024_),
    .Y(_01286_),
    .A1(net278),
    .A2(net781));
 sg13g2_nand2_1 _14317_ (.Y(_08025_),
    .A(\dp.rf.rf[16][9] ),
    .B(net778));
 sg13g2_o21ai_1 _14318_ (.B1(_08025_),
    .Y(_01287_),
    .A1(net273),
    .A2(net778));
 sg13g2_nand2_1 _14319_ (.Y(_08026_),
    .A(\dp.rf.rf[16][10] ),
    .B(net780));
 sg13g2_o21ai_1 _14320_ (.B1(_08026_),
    .Y(_01288_),
    .A1(net270),
    .A2(net780));
 sg13g2_buf_1 fanout250 (.A(net253),
    .X(net250));
 sg13g2_nand2_1 _14322_ (.Y(_08028_),
    .A(\dp.rf.rf[16][11] ),
    .B(net781));
 sg13g2_o21ai_1 _14323_ (.B1(_08028_),
    .Y(_01289_),
    .A1(net263),
    .A2(net781));
 sg13g2_nand2_1 _14324_ (.Y(_08029_),
    .A(\dp.rf.rf[16][12] ),
    .B(net780));
 sg13g2_o21ai_1 _14325_ (.B1(_08029_),
    .Y(_01290_),
    .A1(net256),
    .A2(net780));
 sg13g2_buf_2 fanout249 (.A(net250),
    .X(net249));
 sg13g2_mux2_1 _14327_ (.A0(\dp.rf.rf[16][13] ),
    .A1(net251),
    .S(net773),
    .X(_01291_));
 sg13g2_nor2_1 _14328_ (.A(\dp.rf.rf[16][14] ),
    .B(net772),
    .Y(_08031_));
 sg13g2_a21oi_1 _14329_ (.A1(net246),
    .A2(net772),
    .Y(_01292_),
    .B1(_08031_));
 sg13g2_nand2_1 _14330_ (.Y(_08032_),
    .A(\dp.rf.rf[16][15] ),
    .B(net778));
 sg13g2_o21ai_1 _14331_ (.B1(_08032_),
    .Y(_01293_),
    .A1(net240),
    .A2(net778));
 sg13g2_nand2_1 _14332_ (.Y(_08033_),
    .A(\dp.rf.rf[16][16] ),
    .B(net778));
 sg13g2_o21ai_1 _14333_ (.B1(_08033_),
    .Y(_01294_),
    .A1(net234),
    .A2(net778));
 sg13g2_nand2_1 _14334_ (.Y(_08034_),
    .A(\dp.rf.rf[16][17] ),
    .B(net777));
 sg13g2_o21ai_1 _14335_ (.B1(_08034_),
    .Y(_01295_),
    .A1(net232),
    .A2(net777));
 sg13g2_buf_2 fanout248 (.A(_07550_),
    .X(net248));
 sg13g2_nand2_1 _14337_ (.Y(_08036_),
    .A(\dp.rf.rf[16][18] ),
    .B(net778));
 sg13g2_o21ai_1 _14338_ (.B1(_08036_),
    .Y(_01296_),
    .A1(net227),
    .A2(net778));
 sg13g2_nand2_1 _14339_ (.Y(_08037_),
    .A(\dp.rf.rf[16][19] ),
    .B(net776));
 sg13g2_o21ai_1 _14340_ (.B1(_08037_),
    .Y(_01297_),
    .A1(net222),
    .A2(net776));
 sg13g2_nor2_1 _14341_ (.A(\dp.rf.rf[16][20] ),
    .B(net772),
    .Y(_08038_));
 sg13g2_a21oi_1 _14342_ (.A1(net218),
    .A2(net772),
    .Y(_01298_),
    .B1(_08038_));
 sg13g2_nand2_1 _14343_ (.Y(_08039_),
    .A(\dp.rf.rf[16][21] ),
    .B(net775));
 sg13g2_o21ai_1 _14344_ (.B1(_08039_),
    .Y(_01299_),
    .A1(net211),
    .A2(net775));
 sg13g2_nor2_1 _14345_ (.A(\dp.rf.rf[16][22] ),
    .B(net773),
    .Y(_08040_));
 sg13g2_a21oi_1 _14346_ (.A1(net208),
    .A2(net773),
    .Y(_01300_),
    .B1(_08040_));
 sg13g2_nand2_1 _14347_ (.Y(_08041_),
    .A(\dp.rf.rf[16][23] ),
    .B(net774));
 sg13g2_o21ai_1 _14348_ (.B1(_08041_),
    .Y(_01301_),
    .A1(net203),
    .A2(net774));
 sg13g2_nand2_1 _14349_ (.Y(_08042_),
    .A(\dp.rf.rf[16][24] ),
    .B(net777));
 sg13g2_o21ai_1 _14350_ (.B1(_08042_),
    .Y(_01302_),
    .A1(net197),
    .A2(net777));
 sg13g2_nand2_1 _14351_ (.Y(_08043_),
    .A(\dp.rf.rf[16][25] ),
    .B(net774));
 sg13g2_o21ai_1 _14352_ (.B1(_08043_),
    .Y(_01303_),
    .A1(net190),
    .A2(net774));
 sg13g2_nand2_1 _14353_ (.Y(_08044_),
    .A(\dp.rf.rf[16][26] ),
    .B(net774));
 sg13g2_o21ai_1 _14354_ (.B1(_08044_),
    .Y(_01304_),
    .A1(net185),
    .A2(net774));
 sg13g2_nand2_1 _14355_ (.Y(_08045_),
    .A(\dp.rf.rf[16][27] ),
    .B(net774));
 sg13g2_o21ai_1 _14356_ (.B1(_08045_),
    .Y(_01305_),
    .A1(net180),
    .A2(net774));
 sg13g2_nand2_1 _14357_ (.Y(_08046_),
    .A(\dp.rf.rf[16][28] ),
    .B(net775));
 sg13g2_o21ai_1 _14358_ (.B1(_08046_),
    .Y(_01306_),
    .A1(net308),
    .A2(net775));
 sg13g2_nor2_1 _14359_ (.A(\dp.rf.rf[16][29] ),
    .B(net772),
    .Y(_08047_));
 sg13g2_a21oi_1 _14360_ (.A1(net174),
    .A2(net772),
    .Y(_01307_),
    .B1(_08047_));
 sg13g2_nor2_1 _14361_ (.A(\dp.rf.rf[16][30] ),
    .B(net772),
    .Y(_08048_));
 sg13g2_a21oi_1 _14362_ (.A1(net173),
    .A2(net772),
    .Y(_01308_),
    .B1(_08048_));
 sg13g2_nand2_1 _14363_ (.Y(_08049_),
    .A(\dp.rf.rf[16][31] ),
    .B(net776));
 sg13g2_o21ai_1 _14364_ (.B1(_08049_),
    .Y(_01309_),
    .A1(net167),
    .A2(net776));
 sg13g2_nor2_2 _14365_ (.A(_08015_),
    .B(_07790_),
    .Y(_08050_));
 sg13g2_nor2_1 _14366_ (.A(\dp.rf.rf[17][0] ),
    .B(_08050_),
    .Y(_08051_));
 sg13g2_a21oi_1 _14367_ (.A1(net302),
    .A2(_08050_),
    .Y(_01310_),
    .B1(_08051_));
 sg13g2_nand3_1 _14368_ (.B(_07390_),
    .C(_07789_),
    .A(net1245),
    .Y(_08052_));
 sg13g2_buf_2 fanout247 (.A(net248),
    .X(net247));
 sg13g2_buf_2 fanout246 (.A(_07550_),
    .X(net246));
 sg13g2_buf_2 fanout245 (.A(net246),
    .X(net245));
 sg13g2_nand2_1 _14372_ (.Y(_08056_),
    .A(\dp.rf.rf[17][1] ),
    .B(net770));
 sg13g2_o21ai_1 _14373_ (.B1(_08056_),
    .Y(_01311_),
    .A1(net299),
    .A2(net770));
 sg13g2_nand2_1 _14374_ (.Y(_08057_),
    .A(\dp.rf.rf[17][2] ),
    .B(net771));
 sg13g2_o21ai_1 _14375_ (.B1(_08057_),
    .Y(_01312_),
    .A1(net323),
    .A2(net770));
 sg13g2_nand2_1 _14376_ (.Y(_08058_),
    .A(\dp.rf.rf[17][3] ),
    .B(net770));
 sg13g2_o21ai_1 _14377_ (.B1(_08058_),
    .Y(_01313_),
    .A1(net319),
    .A2(net770));
 sg13g2_and3_1 _14378_ (.X(_08059_),
    .A(net1245),
    .B(_07390_),
    .C(_07789_));
 sg13g2_buf_1 fanout244 (.A(_07558_),
    .X(net244));
 sg13g2_buf_2 fanout243 (.A(net244),
    .X(net243));
 sg13g2_mux2_1 _14381_ (.A0(\dp.rf.rf[17][4] ),
    .A1(net292),
    .S(_08059_),
    .X(_01314_));
 sg13g2_buf_1 fanout242 (.A(_07558_),
    .X(net242));
 sg13g2_nand2_1 _14383_ (.Y(_08063_),
    .A(\dp.rf.rf[17][5] ),
    .B(net768));
 sg13g2_o21ai_1 _14384_ (.B1(_08063_),
    .Y(_01315_),
    .A1(net313),
    .A2(net768));
 sg13g2_nand2_1 _14385_ (.Y(_08064_),
    .A(\dp.rf.rf[17][6] ),
    .B(net768));
 sg13g2_o21ai_1 _14386_ (.B1(_08064_),
    .Y(_01316_),
    .A1(net288),
    .A2(net768));
 sg13g2_nand2_1 _14387_ (.Y(_08065_),
    .A(\dp.rf.rf[17][7] ),
    .B(net769));
 sg13g2_o21ai_1 _14388_ (.B1(_08065_),
    .Y(_01317_),
    .A1(net284),
    .A2(net769));
 sg13g2_nand2_1 _14389_ (.Y(_08066_),
    .A(\dp.rf.rf[17][8] ),
    .B(net770));
 sg13g2_o21ai_1 _14390_ (.B1(_08066_),
    .Y(_01318_),
    .A1(net278),
    .A2(net770));
 sg13g2_nand2_1 _14391_ (.Y(_08067_),
    .A(_07390_),
    .B(_07795_));
 sg13g2_buf_2 fanout241 (.A(net242),
    .X(net241));
 sg13g2_nand2_1 _14393_ (.Y(_08069_),
    .A(\dp.rf.rf[17][9] ),
    .B(net513));
 sg13g2_o21ai_1 _14394_ (.B1(_08069_),
    .Y(_01319_),
    .A1(net271),
    .A2(net513));
 sg13g2_nand2_1 _14395_ (.Y(_08070_),
    .A(\dp.rf.rf[17][10] ),
    .B(net768));
 sg13g2_o21ai_1 _14396_ (.B1(_08070_),
    .Y(_01320_),
    .A1(net268),
    .A2(net768));
 sg13g2_nand2_1 _14397_ (.Y(_08071_),
    .A(\dp.rf.rf[17][11] ),
    .B(net771));
 sg13g2_o21ai_1 _14398_ (.B1(_08071_),
    .Y(_01321_),
    .A1(net263),
    .A2(net770));
 sg13g2_nand2_1 _14399_ (.Y(_08072_),
    .A(\dp.rf.rf[17][12] ),
    .B(net768));
 sg13g2_o21ai_1 _14400_ (.B1(_08072_),
    .Y(_01322_),
    .A1(net257),
    .A2(net768));
 sg13g2_mux2_1 _14401_ (.A0(\dp.rf.rf[17][13] ),
    .A1(net251),
    .S(_08050_),
    .X(_01323_));
 sg13g2_nor2_1 _14402_ (.A(\dp.rf.rf[17][14] ),
    .B(_08050_),
    .Y(_08073_));
 sg13g2_a21oi_1 _14403_ (.A1(net248),
    .A2(_08050_),
    .Y(_01324_),
    .B1(_08073_));
 sg13g2_nand2_1 _14404_ (.Y(_08074_),
    .A(\dp.rf.rf[17][15] ),
    .B(net513));
 sg13g2_o21ai_1 _14405_ (.B1(_08074_),
    .Y(_01325_),
    .A1(net240),
    .A2(net513));
 sg13g2_nand2_1 _14406_ (.Y(_08075_),
    .A(\dp.rf.rf[17][16] ),
    .B(net512));
 sg13g2_o21ai_1 _14407_ (.B1(_08075_),
    .Y(_01326_),
    .A1(net234),
    .A2(net512));
 sg13g2_nor2_1 _14408_ (.A(\dp.rf.rf[17][17] ),
    .B(_08059_),
    .Y(_08076_));
 sg13g2_a21oi_1 _14409_ (.A1(net232),
    .A2(_08059_),
    .Y(_01327_),
    .B1(_08076_));
 sg13g2_nand2_1 _14410_ (.Y(_08077_),
    .A(\dp.rf.rf[17][18] ),
    .B(net769));
 sg13g2_o21ai_1 _14411_ (.B1(_08077_),
    .Y(_01328_),
    .A1(net227),
    .A2(net769));
 sg13g2_nand2_1 _14412_ (.Y(_08078_),
    .A(\dp.rf.rf[17][19] ),
    .B(net767));
 sg13g2_o21ai_1 _14413_ (.B1(_08078_),
    .Y(_01329_),
    .A1(net222),
    .A2(net767));
 sg13g2_nor2_1 _14414_ (.A(\dp.rf.rf[17][20] ),
    .B(net765),
    .Y(_08079_));
 sg13g2_a21oi_1 _14415_ (.A1(net217),
    .A2(net765),
    .Y(_01330_),
    .B1(_08079_));
 sg13g2_nand2_1 _14416_ (.Y(_08080_),
    .A(\dp.rf.rf[17][21] ),
    .B(net766));
 sg13g2_o21ai_1 _14417_ (.B1(_08080_),
    .Y(_01331_),
    .A1(net210),
    .A2(net766));
 sg13g2_nor2_1 _14418_ (.A(\dp.rf.rf[17][22] ),
    .B(net765),
    .Y(_08081_));
 sg13g2_a21oi_1 _14419_ (.A1(net208),
    .A2(net765),
    .Y(_01332_),
    .B1(_08081_));
 sg13g2_nand2_1 _14420_ (.Y(_08082_),
    .A(\dp.rf.rf[17][23] ),
    .B(net512));
 sg13g2_o21ai_1 _14421_ (.B1(_08082_),
    .Y(_01333_),
    .A1(net202),
    .A2(net512));
 sg13g2_nand2_1 _14422_ (.Y(_08083_),
    .A(\dp.rf.rf[17][24] ),
    .B(net767));
 sg13g2_o21ai_1 _14423_ (.B1(_08083_),
    .Y(_01334_),
    .A1(net195),
    .A2(net767));
 sg13g2_nand2_1 _14424_ (.Y(_08084_),
    .A(\dp.rf.rf[17][25] ),
    .B(net766));
 sg13g2_o21ai_1 _14425_ (.B1(_08084_),
    .Y(_01335_),
    .A1(net192),
    .A2(net766));
 sg13g2_nand2_1 _14426_ (.Y(_08085_),
    .A(\dp.rf.rf[17][26] ),
    .B(net512));
 sg13g2_o21ai_1 _14427_ (.B1(_08085_),
    .Y(_01336_),
    .A1(net185),
    .A2(net512));
 sg13g2_nand2_1 _14428_ (.Y(_08086_),
    .A(\dp.rf.rf[17][27] ),
    .B(net766));
 sg13g2_o21ai_1 _14429_ (.B1(_08086_),
    .Y(_01337_),
    .A1(net180),
    .A2(net766));
 sg13g2_nand2_1 _14430_ (.Y(_08087_),
    .A(\dp.rf.rf[17][28] ),
    .B(net766));
 sg13g2_o21ai_1 _14431_ (.B1(_08087_),
    .Y(_01338_),
    .A1(net308),
    .A2(net766));
 sg13g2_nor2_1 _14432_ (.A(\dp.rf.rf[17][29] ),
    .B(net765),
    .Y(_08088_));
 sg13g2_a21oi_1 _14433_ (.A1(net176),
    .A2(net765),
    .Y(_01339_),
    .B1(_08088_));
 sg13g2_nor2_1 _14434_ (.A(\dp.rf.rf[17][30] ),
    .B(net765),
    .Y(_08089_));
 sg13g2_a21oi_1 _14435_ (.A1(net173),
    .A2(net765),
    .Y(_01340_),
    .B1(_08089_));
 sg13g2_nand2_1 _14436_ (.Y(_08090_),
    .A(\dp.rf.rf[17][31] ),
    .B(net512));
 sg13g2_o21ai_1 _14437_ (.B1(_08090_),
    .Y(_01341_),
    .A1(net165),
    .A2(net512));
 sg13g2_nor2_1 _14438_ (.A(_08015_),
    .B(_07924_),
    .Y(_08091_));
 sg13g2_buf_2 fanout240 (.A(net242),
    .X(net240));
 sg13g2_buf_1 fanout239 (.A(_07576_),
    .X(net239));
 sg13g2_nor2_1 _14441_ (.A(\dp.rf.rf[18][0] ),
    .B(_08091_),
    .Y(_08094_));
 sg13g2_a21oi_1 _14442_ (.A1(net302),
    .A2(net511),
    .Y(_01342_),
    .B1(_08094_));
 sg13g2_nand2_1 _14443_ (.Y(_08095_),
    .A(_07390_),
    .B(_07930_));
 sg13g2_buf_1 fanout238 (.A(net239),
    .X(net238));
 sg13g2_buf_2 fanout237 (.A(net239),
    .X(net237));
 sg13g2_buf_2 fanout236 (.A(net238),
    .X(net236));
 sg13g2_nand2_1 _14447_ (.Y(_08099_),
    .A(\dp.rf.rf[18][1] ),
    .B(net763));
 sg13g2_o21ai_1 _14448_ (.B1(_08099_),
    .Y(_01343_),
    .A1(net297),
    .A2(net763));
 sg13g2_nand2_1 _14449_ (.Y(_08100_),
    .A(\dp.rf.rf[18][2] ),
    .B(net764));
 sg13g2_o21ai_1 _14450_ (.B1(_08100_),
    .Y(_01344_),
    .A1(net323),
    .A2(net763));
 sg13g2_nand2_1 _14451_ (.Y(_08101_),
    .A(\dp.rf.rf[18][3] ),
    .B(net763));
 sg13g2_o21ai_1 _14452_ (.B1(_08101_),
    .Y(_01345_),
    .A1(net319),
    .A2(net763));
 sg13g2_mux2_1 _14453_ (.A0(\dp.rf.rf[18][4] ),
    .A1(net290),
    .S(net511),
    .X(_01346_));
 sg13g2_nand2_1 _14454_ (.Y(_08102_),
    .A(\dp.rf.rf[18][5] ),
    .B(net761));
 sg13g2_o21ai_1 _14455_ (.B1(_08102_),
    .Y(_01347_),
    .A1(net314),
    .A2(net761));
 sg13g2_nand2_1 _14456_ (.Y(_08103_),
    .A(\dp.rf.rf[18][6] ),
    .B(net761));
 sg13g2_o21ai_1 _14457_ (.B1(_08103_),
    .Y(_01348_),
    .A1(net288),
    .A2(net761));
 sg13g2_nand2_1 _14458_ (.Y(_08104_),
    .A(\dp.rf.rf[18][7] ),
    .B(net761));
 sg13g2_o21ai_1 _14459_ (.B1(_08104_),
    .Y(_01349_),
    .A1(net284),
    .A2(net761));
 sg13g2_nand2_1 _14460_ (.Y(_08105_),
    .A(\dp.rf.rf[18][8] ),
    .B(net763));
 sg13g2_o21ai_1 _14461_ (.B1(_08105_),
    .Y(_01350_),
    .A1(net279),
    .A2(net763));
 sg13g2_buf_1 fanout235 (.A(net239),
    .X(net235));
 sg13g2_nand2_1 _14463_ (.Y(_08107_),
    .A(\dp.rf.rf[18][9] ),
    .B(net762));
 sg13g2_o21ai_1 _14464_ (.B1(_08107_),
    .Y(_01351_),
    .A1(net271),
    .A2(net762));
 sg13g2_nand2_1 _14465_ (.Y(_08108_),
    .A(\dp.rf.rf[18][10] ),
    .B(net762));
 sg13g2_o21ai_1 _14466_ (.B1(_08108_),
    .Y(_01352_),
    .A1(net270),
    .A2(net764));
 sg13g2_nand2_1 _14467_ (.Y(_08109_),
    .A(\dp.rf.rf[18][11] ),
    .B(net764));
 sg13g2_o21ai_1 _14468_ (.B1(_08109_),
    .Y(_01353_),
    .A1(net263),
    .A2(net763));
 sg13g2_buf_2 fanout234 (.A(net239),
    .X(net234));
 sg13g2_nand2_1 _14470_ (.Y(_08111_),
    .A(\dp.rf.rf[18][12] ),
    .B(net761));
 sg13g2_o21ai_1 _14471_ (.B1(_08111_),
    .Y(_01354_),
    .A1(net257),
    .A2(net761));
 sg13g2_mux2_1 _14472_ (.A0(\dp.rf.rf[18][13] ),
    .A1(net250),
    .S(net511),
    .X(_01355_));
 sg13g2_nor2_1 _14473_ (.A(\dp.rf.rf[18][14] ),
    .B(net510),
    .Y(_08112_));
 sg13g2_a21oi_1 _14474_ (.A1(net246),
    .A2(net510),
    .Y(_01356_),
    .B1(_08112_));
 sg13g2_nand2_1 _14475_ (.Y(_08113_),
    .A(\dp.rf.rf[18][15] ),
    .B(net762));
 sg13g2_o21ai_1 _14476_ (.B1(_08113_),
    .Y(_01357_),
    .A1(net240),
    .A2(net762));
 sg13g2_nand2_1 _14477_ (.Y(_08114_),
    .A(\dp.rf.rf[18][16] ),
    .B(net762));
 sg13g2_o21ai_1 _14478_ (.B1(_08114_),
    .Y(_01358_),
    .A1(net234),
    .A2(net762));
 sg13g2_nor2_1 _14479_ (.A(\dp.rf.rf[18][17] ),
    .B(net511),
    .Y(_08115_));
 sg13g2_a21oi_1 _14480_ (.A1(net232),
    .A2(net511),
    .Y(_01359_),
    .B1(_08115_));
 sg13g2_nand2_1 _14481_ (.Y(_08116_),
    .A(\dp.rf.rf[18][18] ),
    .B(net760));
 sg13g2_o21ai_1 _14482_ (.B1(_08116_),
    .Y(_01360_),
    .A1(net225),
    .A2(net760));
 sg13g2_nand2_1 _14483_ (.Y(_08117_),
    .A(\dp.rf.rf[18][19] ),
    .B(net760));
 sg13g2_o21ai_1 _14484_ (.B1(_08117_),
    .Y(_01361_),
    .A1(net222),
    .A2(net760));
 sg13g2_nor2_1 _14485_ (.A(\dp.rf.rf[18][20] ),
    .B(net510),
    .Y(_08118_));
 sg13g2_a21oi_1 _14486_ (.A1(net217),
    .A2(net510),
    .Y(_01362_),
    .B1(_08118_));
 sg13g2_nand2_1 _14487_ (.Y(_08119_),
    .A(\dp.rf.rf[18][21] ),
    .B(net759));
 sg13g2_o21ai_1 _14488_ (.B1(_08119_),
    .Y(_01363_),
    .A1(net210),
    .A2(net759));
 sg13g2_nor2_1 _14489_ (.A(\dp.rf.rf[18][22] ),
    .B(net510),
    .Y(_08120_));
 sg13g2_a21oi_1 _14490_ (.A1(net208),
    .A2(net511),
    .Y(_01364_),
    .B1(_08120_));
 sg13g2_nand2_1 _14491_ (.Y(_08121_),
    .A(\dp.rf.rf[18][23] ),
    .B(net758));
 sg13g2_o21ai_1 _14492_ (.B1(_08121_),
    .Y(_01365_),
    .A1(net202),
    .A2(net758));
 sg13g2_nand2_1 _14493_ (.Y(_08122_),
    .A(\dp.rf.rf[18][24] ),
    .B(net759));
 sg13g2_o21ai_1 _14494_ (.B1(_08122_),
    .Y(_01366_),
    .A1(net197),
    .A2(net759));
 sg13g2_nand2_1 _14495_ (.Y(_08123_),
    .A(\dp.rf.rf[18][25] ),
    .B(net758));
 sg13g2_o21ai_1 _14496_ (.B1(_08123_),
    .Y(_01367_),
    .A1(net189),
    .A2(net758));
 sg13g2_nand2_1 _14497_ (.Y(_08124_),
    .A(\dp.rf.rf[18][26] ),
    .B(net758));
 sg13g2_o21ai_1 _14498_ (.B1(_08124_),
    .Y(_01368_),
    .A1(net188),
    .A2(net758));
 sg13g2_nand2_1 _14499_ (.Y(_08125_),
    .A(\dp.rf.rf[18][27] ),
    .B(net759));
 sg13g2_o21ai_1 _14500_ (.B1(_08125_),
    .Y(_01369_),
    .A1(net180),
    .A2(net759));
 sg13g2_nand2_1 _14501_ (.Y(_08126_),
    .A(\dp.rf.rf[18][28] ),
    .B(net760));
 sg13g2_o21ai_1 _14502_ (.B1(_08126_),
    .Y(_01370_),
    .A1(net309),
    .A2(net759));
 sg13g2_nor2_1 _14503_ (.A(\dp.rf.rf[18][29] ),
    .B(net510),
    .Y(_08127_));
 sg13g2_a21oi_1 _14504_ (.A1(net176),
    .A2(net511),
    .Y(_01371_),
    .B1(_08127_));
 sg13g2_nor2_1 _14505_ (.A(\dp.rf.rf[18][30] ),
    .B(net510),
    .Y(_08128_));
 sg13g2_a21oi_1 _14506_ (.A1(net172),
    .A2(net510),
    .Y(_01372_),
    .B1(_08128_));
 sg13g2_nand2_1 _14507_ (.Y(_08129_),
    .A(\dp.rf.rf[18][31] ),
    .B(net758));
 sg13g2_o21ai_1 _14508_ (.B1(_08129_),
    .Y(_01373_),
    .A1(net165),
    .A2(net758));
 sg13g2_nand2_1 _14509_ (.Y(_08130_),
    .A(_07795_),
    .B(_07840_));
 sg13g2_buf_1 fanout233 (.A(_07586_),
    .X(net233));
 sg13g2_buf_2 fanout232 (.A(net233),
    .X(net232));
 sg13g2_buf_2 fanout231 (.A(net233),
    .X(net231));
 sg13g2_nand2_1 _14513_ (.Y(_08134_),
    .A(\dp.rf.rf[1][0] ),
    .B(net504));
 sg13g2_o21ai_1 _14514_ (.B1(_08134_),
    .Y(_01374_),
    .A1(net304),
    .A2(net504));
 sg13g2_buf_2 fanout230 (.A(net233),
    .X(net230));
 sg13g2_nand2_1 _14516_ (.Y(_08136_),
    .A(\dp.rf.rf[1][1] ),
    .B(net508));
 sg13g2_o21ai_1 _14517_ (.B1(_08136_),
    .Y(_01375_),
    .A1(net295),
    .A2(net508));
 sg13g2_buf_2 fanout229 (.A(net233),
    .X(net229));
 sg13g2_nand2_1 _14519_ (.Y(_08138_),
    .A(\dp.rf.rf[1][2] ),
    .B(net508));
 sg13g2_o21ai_1 _14520_ (.B1(_08138_),
    .Y(_01376_),
    .A1(net321),
    .A2(net508));
 sg13g2_buf_1 fanout228 (.A(_07599_),
    .X(net228));
 sg13g2_nand2_1 _14522_ (.Y(_08140_),
    .A(\dp.rf.rf[1][3] ),
    .B(net508));
 sg13g2_o21ai_1 _14523_ (.B1(_08140_),
    .Y(_01377_),
    .A1(net315),
    .A2(net508));
 sg13g2_mux2_1 _14524_ (.A0(net294),
    .A1(\dp.rf.rf[1][4] ),
    .S(net507),
    .X(_01378_));
 sg13g2_buf_2 fanout227 (.A(net228),
    .X(net227));
 sg13g2_nand2_1 _14526_ (.Y(_08142_),
    .A(\dp.rf.rf[1][5] ),
    .B(net505));
 sg13g2_o21ai_1 _14527_ (.B1(_08142_),
    .Y(_01379_),
    .A1(net311),
    .A2(net505));
 sg13g2_buf_1 fanout226 (.A(net228),
    .X(net226));
 sg13g2_nand2_1 _14529_ (.Y(_08144_),
    .A(\dp.rf.rf[1][6] ),
    .B(net505));
 sg13g2_o21ai_1 _14530_ (.B1(_08144_),
    .Y(_01380_),
    .A1(net286),
    .A2(net505));
 sg13g2_buf_2 fanout225 (.A(net226),
    .X(net225));
 sg13g2_nand2_1 _14532_ (.Y(_08146_),
    .A(\dp.rf.rf[1][7] ),
    .B(net506));
 sg13g2_o21ai_1 _14533_ (.B1(_08146_),
    .Y(_01381_),
    .A1(net282),
    .A2(net506));
 sg13g2_buf_2 fanout224 (.A(net226),
    .X(net224));
 sg13g2_nand2_1 _14535_ (.Y(_08148_),
    .A(\dp.rf.rf[1][8] ),
    .B(net506));
 sg13g2_o21ai_1 _14536_ (.B1(_08148_),
    .Y(_01382_),
    .A1(net276),
    .A2(net506));
 sg13g2_buf_2 fanout223 (.A(_07608_),
    .X(net223));
 sg13g2_buf_1 fanout222 (.A(net223),
    .X(net222));
 sg13g2_nand2_1 _14539_ (.Y(_08151_),
    .A(\dp.rf.rf[1][9] ),
    .B(net504));
 sg13g2_o21ai_1 _14540_ (.B1(_08151_),
    .Y(_01383_),
    .A1(net274),
    .A2(net504));
 sg13g2_buf_2 fanout221 (.A(net223),
    .X(net221));
 sg13g2_nand2_1 _14542_ (.Y(_08153_),
    .A(\dp.rf.rf[1][10] ),
    .B(net506));
 sg13g2_o21ai_1 _14543_ (.B1(_08153_),
    .Y(_01384_),
    .A1(net266),
    .A2(net506));
 sg13g2_buf_1 fanout220 (.A(_07608_),
    .X(net220));
 sg13g2_buf_2 fanout219 (.A(_07608_),
    .X(net219));
 sg13g2_nand2_1 _14546_ (.Y(_08156_),
    .A(\dp.rf.rf[1][11] ),
    .B(net509));
 sg13g2_o21ai_1 _14547_ (.B1(_08156_),
    .Y(_01385_),
    .A1(net260),
    .A2(net508));
 sg13g2_buf_1 fanout218 (.A(_07620_),
    .X(net218));
 sg13g2_nand2_1 _14549_ (.Y(_08158_),
    .A(\dp.rf.rf[1][12] ),
    .B(net506));
 sg13g2_o21ai_1 _14550_ (.B1(_08158_),
    .Y(_01386_),
    .A1(net254),
    .A2(net506));
 sg13g2_mux2_1 _14551_ (.A0(net252),
    .A1(\dp.rf.rf[1][13] ),
    .S(net508),
    .X(_01387_));
 sg13g2_nand2_1 _14552_ (.Y(_08159_),
    .A(\dp.rf.rf[1][14] ),
    .B(net499));
 sg13g2_o21ai_1 _14553_ (.B1(_08159_),
    .Y(_01388_),
    .A1(net247),
    .A2(net499));
 sg13g2_buf_2 fanout217 (.A(net218),
    .X(net217));
 sg13g2_nand2_1 _14555_ (.Y(_08161_),
    .A(\dp.rf.rf[1][15] ),
    .B(net505));
 sg13g2_o21ai_1 _14556_ (.B1(_08161_),
    .Y(_01389_),
    .A1(net244),
    .A2(net505));
 sg13g2_buf_2 fanout216 (.A(net217),
    .X(net216));
 sg13g2_nand2_1 _14558_ (.Y(_08163_),
    .A(\dp.rf.rf[1][16] ),
    .B(net505));
 sg13g2_o21ai_1 _14559_ (.B1(_08163_),
    .Y(_01390_),
    .A1(net238),
    .A2(net505));
 sg13g2_nand2_1 _14560_ (.Y(_08164_),
    .A(\dp.rf.rf[1][17] ),
    .B(net503));
 sg13g2_o21ai_1 _14561_ (.B1(_08164_),
    .Y(_01391_),
    .A1(net229),
    .A2(net500));
 sg13g2_buf_1 fanout215 (.A(net218),
    .X(net215));
 sg13g2_nand2_1 _14563_ (.Y(_08166_),
    .A(\dp.rf.rf[1][18] ),
    .B(net504));
 sg13g2_o21ai_1 _14564_ (.B1(_08166_),
    .Y(_01392_),
    .A1(net228),
    .A2(net504));
 sg13g2_buf_2 fanout214 (.A(net218),
    .X(net214));
 sg13g2_nand2_1 _14566_ (.Y(_08168_),
    .A(\dp.rf.rf[1][19] ),
    .B(net504));
 sg13g2_o21ai_1 _14567_ (.B1(_08168_),
    .Y(_01393_),
    .A1(net221),
    .A2(net504));
 sg13g2_buf_1 fanout213 (.A(_07630_),
    .X(net213));
 sg13g2_nand2_1 _14569_ (.Y(_08170_),
    .A(\dp.rf.rf[1][20] ),
    .B(net501));
 sg13g2_o21ai_1 _14570_ (.B1(_08170_),
    .Y(_01394_),
    .A1(net215),
    .A2(net501));
 sg13g2_buf_1 fanout212 (.A(net213),
    .X(net212));
 sg13g2_nand2_1 _14572_ (.Y(_08172_),
    .A(\dp.rf.rf[1][21] ),
    .B(net500));
 sg13g2_o21ai_1 _14573_ (.B1(_08172_),
    .Y(_01395_),
    .A1(net213),
    .A2(net500));
 sg13g2_buf_2 fanout211 (.A(net212),
    .X(net211));
 sg13g2_nand2_1 _14575_ (.Y(_08174_),
    .A(\dp.rf.rf[1][22] ),
    .B(net501));
 sg13g2_o21ai_1 _14576_ (.B1(_08174_),
    .Y(_01396_),
    .A1(net206),
    .A2(net502));
 sg13g2_buf_2 fanout210 (.A(net213),
    .X(net210));
 sg13g2_nand2_1 _14578_ (.Y(_08176_),
    .A(\dp.rf.rf[1][23] ),
    .B(net499));
 sg13g2_o21ai_1 _14579_ (.B1(_08176_),
    .Y(_01397_),
    .A1(net203),
    .A2(net499));
 sg13g2_buf_2 fanout209 (.A(net210),
    .X(net209));
 sg13g2_nand2_1 _14581_ (.Y(_08178_),
    .A(\dp.rf.rf[1][24] ),
    .B(net501));
 sg13g2_o21ai_1 _14582_ (.B1(_08178_),
    .Y(_01398_),
    .A1(net196),
    .A2(net501));
 sg13g2_buf_2 fanout208 (.A(_07639_),
    .X(net208));
 sg13g2_nand2_1 _14584_ (.Y(_08180_),
    .A(\dp.rf.rf[1][25] ),
    .B(net500));
 sg13g2_o21ai_1 _14585_ (.B1(_08180_),
    .Y(_01399_),
    .A1(net192),
    .A2(net500));
 sg13g2_buf_2 fanout207 (.A(net208),
    .X(net207));
 sg13g2_nand2_1 _14587_ (.Y(_08182_),
    .A(\dp.rf.rf[1][26] ),
    .B(net501));
 sg13g2_o21ai_1 _14588_ (.B1(_08182_),
    .Y(_01400_),
    .A1(net186),
    .A2(net501));
 sg13g2_buf_2 fanout206 (.A(_07639_),
    .X(net206));
 sg13g2_nand2_1 _14590_ (.Y(_08184_),
    .A(\dp.rf.rf[1][27] ),
    .B(net499));
 sg13g2_o21ai_1 _14591_ (.B1(_08184_),
    .Y(_01401_),
    .A1(net181),
    .A2(net499));
 sg13g2_buf_2 fanout205 (.A(net206),
    .X(net205));
 sg13g2_nand2_1 _14593_ (.Y(_08186_),
    .A(\dp.rf.rf[1][28] ),
    .B(net500));
 sg13g2_o21ai_1 _14594_ (.B1(_08186_),
    .Y(_01402_),
    .A1(net307),
    .A2(net500));
 sg13g2_nand2_1 _14595_ (.Y(_08187_),
    .A(\dp.rf.rf[1][29] ),
    .B(net502));
 sg13g2_o21ai_1 _14596_ (.B1(_08187_),
    .Y(_01403_),
    .A1(net177),
    .A2(net502));
 sg13g2_nand2_1 _14597_ (.Y(_08188_),
    .A(\dp.rf.rf[1][30] ),
    .B(net501));
 sg13g2_o21ai_1 _14598_ (.B1(_08188_),
    .Y(_01404_),
    .A1(net171),
    .A2(net502));
 sg13g2_buf_1 fanout204 (.A(_07650_),
    .X(net204));
 sg13g2_nand2_1 _14600_ (.Y(_08190_),
    .A(\dp.rf.rf[1][31] ),
    .B(net499));
 sg13g2_o21ai_1 _14601_ (.B1(_08190_),
    .Y(_01405_),
    .A1(net168),
    .A2(net499));
 sg13g2_nor3_2 _14602_ (.A(_05285_),
    .B(net1256),
    .C(_05508_),
    .Y(_08191_));
 sg13g2_nand2_1 _14603_ (.Y(_08192_),
    .A(_07841_),
    .B(_08191_));
 sg13g2_buf_2 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_2 fanout202 (.A(net204),
    .X(net202));
 sg13g2_buf_1 fanout201 (.A(_07650_),
    .X(net201));
 sg13g2_nand2_1 _14607_ (.Y(_08196_),
    .A(\dp.rf.rf[20][0] ),
    .B(net754));
 sg13g2_o21ai_1 _14608_ (.B1(_08196_),
    .Y(_01406_),
    .A1(net301),
    .A2(net754));
 sg13g2_nand2_1 _14609_ (.Y(_08197_),
    .A(\dp.rf.rf[20][1] ),
    .B(net755));
 sg13g2_o21ai_1 _14610_ (.B1(_08197_),
    .Y(_01407_),
    .A1(net297),
    .A2(net755));
 sg13g2_buf_2 fanout200 (.A(_07650_),
    .X(net200));
 sg13g2_nand2_1 _14612_ (.Y(_08199_),
    .A(\dp.rf.rf[20][2] ),
    .B(net756));
 sg13g2_o21ai_1 _14613_ (.B1(_08199_),
    .Y(_01408_),
    .A1(net323),
    .A2(net755));
 sg13g2_nand2_1 _14614_ (.Y(_08200_),
    .A(\dp.rf.rf[20][3] ),
    .B(net755));
 sg13g2_o21ai_1 _14615_ (.B1(_08200_),
    .Y(_01409_),
    .A1(net319),
    .A2(net755));
 sg13g2_nand3b_1 _14616_ (.B(net1244),
    .C(net1247),
    .Y(_08201_),
    .A_N(net1256));
 sg13g2_buf_1 fanout199 (.A(_07660_),
    .X(net199));
 sg13g2_nor2_2 _14618_ (.A(_08016_),
    .B(_08201_),
    .Y(_08203_));
 sg13g2_buf_2 fanout198 (.A(net199),
    .X(net198));
 sg13g2_mux2_1 _14620_ (.A0(\dp.rf.rf[20][4] ),
    .A1(net291),
    .S(_08203_),
    .X(_01410_));
 sg13g2_nand2_1 _14621_ (.Y(_08205_),
    .A(\dp.rf.rf[20][5] ),
    .B(net753));
 sg13g2_o21ai_1 _14622_ (.B1(_08205_),
    .Y(_01411_),
    .A1(net313),
    .A2(net753));
 sg13g2_nand2_1 _14623_ (.Y(_08206_),
    .A(\dp.rf.rf[20][6] ),
    .B(net753));
 sg13g2_o21ai_1 _14624_ (.B1(_08206_),
    .Y(_01412_),
    .A1(net287),
    .A2(net753));
 sg13g2_nand2_1 _14625_ (.Y(_08207_),
    .A(\dp.rf.rf[20][7] ),
    .B(net754));
 sg13g2_o21ai_1 _14626_ (.B1(_08207_),
    .Y(_01413_),
    .A1(net283),
    .A2(net757));
 sg13g2_nand2_1 _14627_ (.Y(_08208_),
    .A(\dp.rf.rf[20][8] ),
    .B(net756));
 sg13g2_o21ai_1 _14628_ (.B1(_08208_),
    .Y(_01414_),
    .A1(net277),
    .A2(net756));
 sg13g2_nand2_1 _14629_ (.Y(_08209_),
    .A(\dp.rf.rf[20][9] ),
    .B(net754));
 sg13g2_o21ai_1 _14630_ (.B1(_08209_),
    .Y(_01415_),
    .A1(net272),
    .A2(net754));
 sg13g2_nand2_1 _14631_ (.Y(_08210_),
    .A(\dp.rf.rf[20][10] ),
    .B(net755));
 sg13g2_o21ai_1 _14632_ (.B1(_08210_),
    .Y(_01416_),
    .A1(net269),
    .A2(net755));
 sg13g2_buf_2 fanout197 (.A(net198),
    .X(net197));
 sg13g2_nand2_1 _14634_ (.Y(_08212_),
    .A(\dp.rf.rf[20][11] ),
    .B(net755));
 sg13g2_o21ai_1 _14635_ (.B1(_08212_),
    .Y(_01417_),
    .A1(net264),
    .A2(net756));
 sg13g2_nand2_1 _14636_ (.Y(_08213_),
    .A(\dp.rf.rf[20][12] ),
    .B(net753));
 sg13g2_o21ai_1 _14637_ (.B1(_08213_),
    .Y(_01418_),
    .A1(net258),
    .A2(net753));
 sg13g2_mux2_1 _14638_ (.A0(\dp.rf.rf[20][13] ),
    .A1(net253),
    .S(_08203_),
    .X(_01419_));
 sg13g2_buf_2 fanout196 (.A(net199),
    .X(net196));
 sg13g2_nand2_1 _14640_ (.Y(_08215_),
    .A(\dp.rf.rf[20][14] ),
    .B(net750));
 sg13g2_o21ai_1 _14641_ (.B1(_08215_),
    .Y(_01420_),
    .A1(net245),
    .A2(net750));
 sg13g2_nand2_1 _14642_ (.Y(_08216_),
    .A(\dp.rf.rf[20][15] ),
    .B(net753));
 sg13g2_o21ai_1 _14643_ (.B1(_08216_),
    .Y(_01421_),
    .A1(net240),
    .A2(net753));
 sg13g2_nand2_1 _14644_ (.Y(_08217_),
    .A(\dp.rf.rf[20][16] ),
    .B(net754));
 sg13g2_o21ai_1 _14645_ (.B1(_08217_),
    .Y(_01422_),
    .A1(net237),
    .A2(net754));
 sg13g2_nand2_1 _14646_ (.Y(_08218_),
    .A(\dp.rf.rf[20][17] ),
    .B(net752));
 sg13g2_o21ai_1 _14647_ (.B1(_08218_),
    .Y(_01423_),
    .A1(net229),
    .A2(net752));
 sg13g2_nand2_1 _14648_ (.Y(_08219_),
    .A(\dp.rf.rf[20][18] ),
    .B(net751));
 sg13g2_o21ai_1 _14649_ (.B1(_08219_),
    .Y(_01424_),
    .A1(net224),
    .A2(net751));
 sg13g2_nand2_1 _14650_ (.Y(_08220_),
    .A(\dp.rf.rf[20][19] ),
    .B(net751));
 sg13g2_o21ai_1 _14651_ (.B1(_08220_),
    .Y(_01425_),
    .A1(net221),
    .A2(net751));
 sg13g2_nand2_1 _14652_ (.Y(_08221_),
    .A(\dp.rf.rf[20][20] ),
    .B(net757));
 sg13g2_o21ai_1 _14653_ (.B1(_08221_),
    .Y(_01426_),
    .A1(net216),
    .A2(net752));
 sg13g2_nand2_1 _14654_ (.Y(_08222_),
    .A(\dp.rf.rf[20][21] ),
    .B(net750));
 sg13g2_o21ai_1 _14655_ (.B1(_08222_),
    .Y(_01427_),
    .A1(net211),
    .A2(net750));
 sg13g2_nor2_1 _14656_ (.A(\dp.rf.rf[20][22] ),
    .B(_08203_),
    .Y(_08223_));
 sg13g2_a21oi_1 _14657_ (.A1(net208),
    .A2(_08203_),
    .Y(_01428_),
    .B1(_08223_));
 sg13g2_nand2_1 _14658_ (.Y(_08224_),
    .A(\dp.rf.rf[20][23] ),
    .B(net749));
 sg13g2_o21ai_1 _14659_ (.B1(_08224_),
    .Y(_01429_),
    .A1(net200),
    .A2(net749));
 sg13g2_nand2_1 _14660_ (.Y(_08225_),
    .A(\dp.rf.rf[20][24] ),
    .B(net752));
 sg13g2_o21ai_1 _14661_ (.B1(_08225_),
    .Y(_01430_),
    .A1(net198),
    .A2(net752));
 sg13g2_nand2_1 _14662_ (.Y(_08226_),
    .A(\dp.rf.rf[20][25] ),
    .B(net749));
 sg13g2_o21ai_1 _14663_ (.B1(_08226_),
    .Y(_01431_),
    .A1(net189),
    .A2(net749));
 sg13g2_nand2_1 _14664_ (.Y(_08227_),
    .A(\dp.rf.rf[20][26] ),
    .B(net749));
 sg13g2_o21ai_1 _14665_ (.B1(_08227_),
    .Y(_01432_),
    .A1(net183),
    .A2(net749));
 sg13g2_nand2_1 _14666_ (.Y(_08228_),
    .A(\dp.rf.rf[20][27] ),
    .B(net749));
 sg13g2_o21ai_1 _14667_ (.B1(_08228_),
    .Y(_01433_),
    .A1(net179),
    .A2(net749));
 sg13g2_nand2_1 _14668_ (.Y(_08229_),
    .A(\dp.rf.rf[20][28] ),
    .B(net750));
 sg13g2_o21ai_1 _14669_ (.B1(_08229_),
    .Y(_01434_),
    .A1(net306),
    .A2(net750));
 sg13g2_nor2_1 _14670_ (.A(\dp.rf.rf[20][29] ),
    .B(_08203_),
    .Y(_08230_));
 sg13g2_a21oi_1 _14671_ (.A1(net174),
    .A2(_08203_),
    .Y(_01435_),
    .B1(_08230_));
 sg13g2_nand2_1 _14672_ (.Y(_08231_),
    .A(\dp.rf.rf[20][30] ),
    .B(net752));
 sg13g2_o21ai_1 _14673_ (.B1(_08231_),
    .Y(_01436_),
    .A1(net172),
    .A2(net752));
 sg13g2_nand2_1 _14674_ (.Y(_08232_),
    .A(\dp.rf.rf[20][31] ),
    .B(net751));
 sg13g2_o21ai_1 _14675_ (.B1(_08232_),
    .Y(_01437_),
    .A1(net165),
    .A2(net751));
 sg13g2_nand2_1 _14676_ (.Y(_08233_),
    .A(_07746_),
    .B(_07841_));
 sg13g2_buf_2 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_1 fanout194 (.A(_07677_),
    .X(net194));
 sg13g2_buf_1 fanout193 (.A(net194),
    .X(net193));
 sg13g2_nand2_1 _14680_ (.Y(_08237_),
    .A(\dp.rf.rf[8][0] ),
    .B(net746));
 sg13g2_o21ai_1 _14681_ (.B1(_08237_),
    .Y(_01438_),
    .A1(net300),
    .A2(net746));
 sg13g2_nand2_1 _14682_ (.Y(_08238_),
    .A(\dp.rf.rf[8][1] ),
    .B(net748));
 sg13g2_o21ai_1 _14683_ (.B1(_08238_),
    .Y(_01439_),
    .A1(net295),
    .A2(net747));
 sg13g2_nand2_1 _14684_ (.Y(_08239_),
    .A(\dp.rf.rf[8][2] ),
    .B(net748));
 sg13g2_o21ai_1 _14685_ (.B1(_08239_),
    .Y(_01440_),
    .A1(net320),
    .A2(net747));
 sg13g2_nand2_1 _14686_ (.Y(_08240_),
    .A(\dp.rf.rf[8][3] ),
    .B(net747));
 sg13g2_o21ai_1 _14687_ (.B1(_08240_),
    .Y(_01441_),
    .A1(net315),
    .A2(net747));
 sg13g2_mux2_1 _14688_ (.A0(net294),
    .A1(\dp.rf.rf[8][4] ),
    .S(net746),
    .X(_01442_));
 sg13g2_nand2_1 _14689_ (.Y(_08241_),
    .A(\dp.rf.rf[8][5] ),
    .B(net743));
 sg13g2_o21ai_1 _14690_ (.B1(_08241_),
    .Y(_01443_),
    .A1(net310),
    .A2(net744));
 sg13g2_nand2_1 _14691_ (.Y(_08242_),
    .A(\dp.rf.rf[8][6] ),
    .B(net744));
 sg13g2_o21ai_1 _14692_ (.B1(_08242_),
    .Y(_01444_),
    .A1(net286),
    .A2(net743));
 sg13g2_nand2_1 _14693_ (.Y(_08243_),
    .A(\dp.rf.rf[8][7] ),
    .B(net743));
 sg13g2_o21ai_1 _14694_ (.B1(_08243_),
    .Y(_01445_),
    .A1(net281),
    .A2(net743));
 sg13g2_nand2_1 _14695_ (.Y(_08244_),
    .A(\dp.rf.rf[8][8] ),
    .B(net745));
 sg13g2_o21ai_1 _14696_ (.B1(_08244_),
    .Y(_01446_),
    .A1(net276),
    .A2(net745));
 sg13g2_buf_2 fanout192 (.A(net193),
    .X(net192));
 sg13g2_nand2_1 _14698_ (.Y(_08246_),
    .A(\dp.rf.rf[8][9] ),
    .B(net743));
 sg13g2_o21ai_1 _14699_ (.B1(_08246_),
    .Y(_01447_),
    .A1(net274),
    .A2(net743));
 sg13g2_nand2_1 _14700_ (.Y(_08247_),
    .A(\dp.rf.rf[8][10] ),
    .B(net745));
 sg13g2_o21ai_1 _14701_ (.B1(_08247_),
    .Y(_01448_),
    .A1(net266),
    .A2(net745));
 sg13g2_buf_2 fanout191 (.A(net194),
    .X(net191));
 sg13g2_nand2_1 _14703_ (.Y(_08249_),
    .A(\dp.rf.rf[8][11] ),
    .B(net747));
 sg13g2_o21ai_1 _14704_ (.B1(_08249_),
    .Y(_01449_),
    .A1(net260),
    .A2(net747));
 sg13g2_nand2_1 _14705_ (.Y(_08250_),
    .A(\dp.rf.rf[8][12] ),
    .B(net745));
 sg13g2_o21ai_1 _14706_ (.B1(_08250_),
    .Y(_01450_),
    .A1(net254),
    .A2(net745));
 sg13g2_mux2_1 _14707_ (.A0(net249),
    .A1(\dp.rf.rf[8][13] ),
    .S(net746),
    .X(_01451_));
 sg13g2_nand2_1 _14708_ (.Y(_08251_),
    .A(\dp.rf.rf[8][14] ),
    .B(net740));
 sg13g2_o21ai_1 _14709_ (.B1(_08251_),
    .Y(_01452_),
    .A1(net247),
    .A2(net740));
 sg13g2_nand2_1 _14710_ (.Y(_08252_),
    .A(\dp.rf.rf[8][15] ),
    .B(net744));
 sg13g2_o21ai_1 _14711_ (.B1(_08252_),
    .Y(_01453_),
    .A1(net244),
    .A2(net744));
 sg13g2_nand2_1 _14712_ (.Y(_08253_),
    .A(\dp.rf.rf[8][16] ),
    .B(net743));
 sg13g2_o21ai_1 _14713_ (.B1(_08253_),
    .Y(_01454_),
    .A1(net237),
    .A2(net743));
 sg13g2_nand2_1 _14714_ (.Y(_08254_),
    .A(\dp.rf.rf[8][17] ),
    .B(net742));
 sg13g2_o21ai_1 _14715_ (.B1(_08254_),
    .Y(_01455_),
    .A1(net229),
    .A2(net742));
 sg13g2_nand2_1 _14716_ (.Y(_08255_),
    .A(\dp.rf.rf[8][18] ),
    .B(net746));
 sg13g2_o21ai_1 _14717_ (.B1(_08255_),
    .Y(_01456_),
    .A1(net227),
    .A2(net746));
 sg13g2_nand2_1 _14718_ (.Y(_08256_),
    .A(\dp.rf.rf[8][19] ),
    .B(net746));
 sg13g2_o21ai_1 _14719_ (.B1(_08256_),
    .Y(_01457_),
    .A1(net219),
    .A2(net746));
 sg13g2_buf_1 fanout190 (.A(net194),
    .X(net190));
 sg13g2_nand2_1 _14721_ (.Y(_08258_),
    .A(\dp.rf.rf[8][20] ),
    .B(net741));
 sg13g2_o21ai_1 _14722_ (.B1(_08258_),
    .Y(_01458_),
    .A1(net214),
    .A2(net741));
 sg13g2_nand2_1 _14723_ (.Y(_08259_),
    .A(\dp.rf.rf[8][21] ),
    .B(net739));
 sg13g2_o21ai_1 _14724_ (.B1(_08259_),
    .Y(_01459_),
    .A1(net209),
    .A2(net739));
 sg13g2_buf_2 fanout189 (.A(net194),
    .X(net189));
 sg13g2_nand2_1 _14726_ (.Y(_08261_),
    .A(\dp.rf.rf[8][22] ),
    .B(net741));
 sg13g2_o21ai_1 _14727_ (.B1(_08261_),
    .Y(_01460_),
    .A1(net205),
    .A2(net742));
 sg13g2_nand2_1 _14728_ (.Y(_08262_),
    .A(\dp.rf.rf[8][23] ),
    .B(net740));
 sg13g2_o21ai_1 _14729_ (.B1(_08262_),
    .Y(_01461_),
    .A1(net204),
    .A2(net740));
 sg13g2_nand2_1 _14730_ (.Y(_08263_),
    .A(\dp.rf.rf[8][24] ),
    .B(net739));
 sg13g2_o21ai_1 _14731_ (.B1(_08263_),
    .Y(_01462_),
    .A1(net199),
    .A2(net739));
 sg13g2_nand2_1 _14732_ (.Y(_08264_),
    .A(\dp.rf.rf[8][25] ),
    .B(net739));
 sg13g2_o21ai_1 _14733_ (.B1(_08264_),
    .Y(_01463_),
    .A1(net192),
    .A2(net739));
 sg13g2_nand2_1 _14734_ (.Y(_08265_),
    .A(\dp.rf.rf[8][26] ),
    .B(net741));
 sg13g2_o21ai_1 _14735_ (.B1(_08265_),
    .Y(_01464_),
    .A1(net187),
    .A2(net741));
 sg13g2_nand2_1 _14736_ (.Y(_08266_),
    .A(\dp.rf.rf[8][27] ),
    .B(net740));
 sg13g2_o21ai_1 _14737_ (.B1(_08266_),
    .Y(_01465_),
    .A1(net181),
    .A2(net740));
 sg13g2_nand2_1 _14738_ (.Y(_08267_),
    .A(\dp.rf.rf[8][28] ),
    .B(net739));
 sg13g2_o21ai_1 _14739_ (.B1(_08267_),
    .Y(_01466_),
    .A1(net309),
    .A2(net739));
 sg13g2_nand2_1 _14740_ (.Y(_08268_),
    .A(\dp.rf.rf[8][29] ),
    .B(net741));
 sg13g2_o21ai_1 _14741_ (.B1(_08268_),
    .Y(_01467_),
    .A1(net178),
    .A2(net742));
 sg13g2_nand2_1 _14742_ (.Y(_08269_),
    .A(\dp.rf.rf[8][30] ),
    .B(net741));
 sg13g2_o21ai_1 _14743_ (.B1(_08269_),
    .Y(_01468_),
    .A1(net170),
    .A2(net741));
 sg13g2_nand2_1 _14744_ (.Y(_08270_),
    .A(\dp.rf.rf[8][31] ),
    .B(net740));
 sg13g2_o21ai_1 _14745_ (.B1(_08270_),
    .Y(_01469_),
    .A1(net168),
    .A2(net740));
 sg13g2_nand2_1 _14746_ (.Y(_08271_),
    .A(_07746_),
    .B(_07930_));
 sg13g2_buf_1 fanout188 (.A(_07686_),
    .X(net188));
 sg13g2_buf_2 fanout187 (.A(net188),
    .X(net187));
 sg13g2_buf_2 fanout186 (.A(net187),
    .X(net186));
 sg13g2_nand2_1 _14750_ (.Y(_08275_),
    .A(\dp.rf.rf[10][0] ),
    .B(net736));
 sg13g2_o21ai_1 _14751_ (.B1(_08275_),
    .Y(_01470_),
    .A1(net300),
    .A2(net736));
 sg13g2_nand2_1 _14752_ (.Y(_08276_),
    .A(\dp.rf.rf[10][1] ),
    .B(net737));
 sg13g2_o21ai_1 _14753_ (.B1(_08276_),
    .Y(_01471_),
    .A1(net295),
    .A2(net737));
 sg13g2_nand2_1 _14754_ (.Y(_08277_),
    .A(\dp.rf.rf[10][2] ),
    .B(net737));
 sg13g2_o21ai_1 _14755_ (.B1(_08277_),
    .Y(_01472_),
    .A1(net320),
    .A2(net737));
 sg13g2_nand2_1 _14756_ (.Y(_08278_),
    .A(\dp.rf.rf[10][3] ),
    .B(net738));
 sg13g2_o21ai_1 _14757_ (.B1(_08278_),
    .Y(_01473_),
    .A1(net315),
    .A2(net738));
 sg13g2_mux2_1 _14758_ (.A0(net294),
    .A1(\dp.rf.rf[10][4] ),
    .S(net736),
    .X(_01474_));
 sg13g2_nand2_1 _14759_ (.Y(_08279_),
    .A(\dp.rf.rf[10][5] ),
    .B(net734));
 sg13g2_o21ai_1 _14760_ (.B1(_08279_),
    .Y(_01475_),
    .A1(net310),
    .A2(net734));
 sg13g2_nand2_1 _14761_ (.Y(_08280_),
    .A(\dp.rf.rf[10][6] ),
    .B(net733));
 sg13g2_o21ai_1 _14762_ (.B1(_08280_),
    .Y(_01476_),
    .A1(net286),
    .A2(net733));
 sg13g2_nand2_1 _14763_ (.Y(_08281_),
    .A(\dp.rf.rf[10][7] ),
    .B(net733));
 sg13g2_o21ai_1 _14764_ (.B1(_08281_),
    .Y(_01477_),
    .A1(net281),
    .A2(net733));
 sg13g2_nand2_1 _14765_ (.Y(_08282_),
    .A(\dp.rf.rf[10][8] ),
    .B(net735));
 sg13g2_o21ai_1 _14766_ (.B1(_08282_),
    .Y(_01478_),
    .A1(net276),
    .A2(net735));
 sg13g2_buf_1 fanout185 (.A(net188),
    .X(net185));
 sg13g2_nand2_1 _14768_ (.Y(_08284_),
    .A(\dp.rf.rf[10][9] ),
    .B(net733));
 sg13g2_o21ai_1 _14769_ (.B1(_08284_),
    .Y(_01479_),
    .A1(net274),
    .A2(net733));
 sg13g2_nand2_1 _14770_ (.Y(_08285_),
    .A(\dp.rf.rf[10][10] ),
    .B(net735));
 sg13g2_o21ai_1 _14771_ (.B1(_08285_),
    .Y(_01480_),
    .A1(net266),
    .A2(net735));
 sg13g2_buf_1 fanout184 (.A(net185),
    .X(net184));
 sg13g2_nand2_1 _14773_ (.Y(_08287_),
    .A(\dp.rf.rf[10][11] ),
    .B(net737));
 sg13g2_o21ai_1 _14774_ (.B1(_08287_),
    .Y(_01481_),
    .A1(net260),
    .A2(net737));
 sg13g2_nand2_1 _14775_ (.Y(_08288_),
    .A(\dp.rf.rf[10][12] ),
    .B(net737));
 sg13g2_o21ai_1 _14776_ (.B1(_08288_),
    .Y(_01482_),
    .A1(net254),
    .A2(net737));
 sg13g2_mux2_1 _14777_ (.A0(net249),
    .A1(\dp.rf.rf[10][13] ),
    .S(net736),
    .X(_01483_));
 sg13g2_nand2_1 _14778_ (.Y(_08289_),
    .A(\dp.rf.rf[10][14] ),
    .B(net728));
 sg13g2_o21ai_1 _14779_ (.B1(_08289_),
    .Y(_01484_),
    .A1(net248),
    .A2(net728));
 sg13g2_nand2_1 _14780_ (.Y(_08290_),
    .A(\dp.rf.rf[10][15] ),
    .B(net734));
 sg13g2_o21ai_1 _14781_ (.B1(_08290_),
    .Y(_01485_),
    .A1(net243),
    .A2(net734));
 sg13g2_nand2_1 _14782_ (.Y(_08291_),
    .A(\dp.rf.rf[10][16] ),
    .B(net733));
 sg13g2_o21ai_1 _14783_ (.B1(_08291_),
    .Y(_01486_),
    .A1(net237),
    .A2(net733));
 sg13g2_nand2_1 _14784_ (.Y(_08292_),
    .A(\dp.rf.rf[10][17] ),
    .B(net729));
 sg13g2_o21ai_1 _14785_ (.B1(_08292_),
    .Y(_01487_),
    .A1(net229),
    .A2(net729));
 sg13g2_nand2_1 _14786_ (.Y(_08293_),
    .A(\dp.rf.rf[10][18] ),
    .B(net736));
 sg13g2_o21ai_1 _14787_ (.B1(_08293_),
    .Y(_01488_),
    .A1(net227),
    .A2(net736));
 sg13g2_nand2_1 _14788_ (.Y(_08294_),
    .A(\dp.rf.rf[10][19] ),
    .B(net736));
 sg13g2_o21ai_1 _14789_ (.B1(_08294_),
    .Y(_01489_),
    .A1(net219),
    .A2(net736));
 sg13g2_buf_2 fanout183 (.A(net185),
    .X(net183));
 sg13g2_nand2_1 _14791_ (.Y(_08296_),
    .A(\dp.rf.rf[10][20] ),
    .B(net731));
 sg13g2_o21ai_1 _14792_ (.B1(_08296_),
    .Y(_01490_),
    .A1(net214),
    .A2(net731));
 sg13g2_nand2_1 _14793_ (.Y(_08297_),
    .A(\dp.rf.rf[10][21] ),
    .B(net730));
 sg13g2_o21ai_1 _14794_ (.B1(_08297_),
    .Y(_01491_),
    .A1(net209),
    .A2(net730));
 sg13g2_buf_2 fanout182 (.A(_07697_),
    .X(net182));
 sg13g2_buf_2 fanout181 (.A(net182),
    .X(net181));
 sg13g2_nand2_1 _14797_ (.Y(_08300_),
    .A(\dp.rf.rf[10][22] ),
    .B(net732));
 sg13g2_o21ai_1 _14798_ (.B1(_08300_),
    .Y(_01492_),
    .A1(net205),
    .A2(net732));
 sg13g2_nand2_1 _14799_ (.Y(_08301_),
    .A(\dp.rf.rf[10][23] ),
    .B(net728));
 sg13g2_o21ai_1 _14800_ (.B1(_08301_),
    .Y(_01493_),
    .A1(net203),
    .A2(net728));
 sg13g2_nand2_1 _14801_ (.Y(_08302_),
    .A(\dp.rf.rf[10][24] ),
    .B(net730));
 sg13g2_o21ai_1 _14802_ (.B1(_08302_),
    .Y(_01494_),
    .A1(net196),
    .A2(net730));
 sg13g2_nand2_1 _14803_ (.Y(_08303_),
    .A(\dp.rf.rf[10][25] ),
    .B(net730));
 sg13g2_o21ai_1 _14804_ (.B1(_08303_),
    .Y(_01495_),
    .A1(net193),
    .A2(net730));
 sg13g2_nand2_1 _14805_ (.Y(_08304_),
    .A(\dp.rf.rf[10][26] ),
    .B(net731));
 sg13g2_o21ai_1 _14806_ (.B1(_08304_),
    .Y(_01496_),
    .A1(net186),
    .A2(net731));
 sg13g2_nand2_1 _14807_ (.Y(_08305_),
    .A(\dp.rf.rf[10][27] ),
    .B(net728));
 sg13g2_o21ai_1 _14808_ (.B1(_08305_),
    .Y(_01497_),
    .A1(net181),
    .A2(net728));
 sg13g2_nand2_1 _14809_ (.Y(_08306_),
    .A(\dp.rf.rf[10][28] ),
    .B(net729));
 sg13g2_o21ai_1 _14810_ (.B1(_08306_),
    .Y(_01498_),
    .A1(net307),
    .A2(net729));
 sg13g2_buf_2 fanout180 (.A(_07697_),
    .X(net180));
 sg13g2_nand2_1 _14812_ (.Y(_08308_),
    .A(\dp.rf.rf[10][29] ),
    .B(net731));
 sg13g2_o21ai_1 _14813_ (.B1(_08308_),
    .Y(_01499_),
    .A1(net178),
    .A2(net731));
 sg13g2_nand2_1 _14814_ (.Y(_08309_),
    .A(\dp.rf.rf[10][30] ),
    .B(net731));
 sg13g2_o21ai_1 _14815_ (.B1(_08309_),
    .Y(_01500_),
    .A1(net170),
    .A2(net731));
 sg13g2_nand2_1 _14816_ (.Y(_08310_),
    .A(\dp.rf.rf[10][31] ),
    .B(net728));
 sg13g2_o21ai_1 _14817_ (.B1(_08310_),
    .Y(_01501_),
    .A1(net168),
    .A2(net728));
 sg13g2_nor3_2 _14818_ (.A(net1247),
    .B(net1257),
    .C(_05508_),
    .Y(_08311_));
 sg13g2_nand2_1 _14819_ (.Y(_08312_),
    .A(_07396_),
    .B(_08311_));
 sg13g2_buf_2 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_2 fanout178 (.A(_07719_),
    .X(net178));
 sg13g2_buf_2 fanout177 (.A(net178),
    .X(net177));
 sg13g2_nand2_1 _14823_ (.Y(_08316_),
    .A(\dp.rf.rf[7][0] ),
    .B(net495));
 sg13g2_o21ai_1 _14824_ (.B1(_08316_),
    .Y(_01502_),
    .A1(net303),
    .A2(net495));
 sg13g2_nand2_1 _14825_ (.Y(_08317_),
    .A(\dp.rf.rf[7][1] ),
    .B(net496));
 sg13g2_o21ai_1 _14826_ (.B1(_08317_),
    .Y(_01503_),
    .A1(net296),
    .A2(net496));
 sg13g2_nand2_1 _14827_ (.Y(_08318_),
    .A(\dp.rf.rf[7][2] ),
    .B(net496));
 sg13g2_o21ai_1 _14828_ (.B1(_08318_),
    .Y(_01504_),
    .A1(net320),
    .A2(net496));
 sg13g2_nand2_1 _14829_ (.Y(_08319_),
    .A(\dp.rf.rf[7][3] ),
    .B(net497));
 sg13g2_o21ai_1 _14830_ (.B1(_08319_),
    .Y(_01505_),
    .A1(net316),
    .A2(net496));
 sg13g2_mux2_1 _14831_ (.A0(net290),
    .A1(\dp.rf.rf[7][4] ),
    .S(net490),
    .X(_01506_));
 sg13g2_nand2_1 _14832_ (.Y(_08320_),
    .A(\dp.rf.rf[7][5] ),
    .B(net494));
 sg13g2_o21ai_1 _14833_ (.B1(_08320_),
    .Y(_01507_),
    .A1(net311),
    .A2(net494));
 sg13g2_nand2_1 _14834_ (.Y(_08321_),
    .A(\dp.rf.rf[7][6] ),
    .B(net493));
 sg13g2_o21ai_1 _14835_ (.B1(_08321_),
    .Y(_01508_),
    .A1(net285),
    .A2(net493));
 sg13g2_nand2_1 _14836_ (.Y(_08322_),
    .A(\dp.rf.rf[7][7] ),
    .B(net493));
 sg13g2_o21ai_1 _14837_ (.B1(_08322_),
    .Y(_01509_),
    .A1(net282),
    .A2(net493));
 sg13g2_nand2_1 _14838_ (.Y(_08323_),
    .A(\dp.rf.rf[7][8] ),
    .B(net496));
 sg13g2_o21ai_1 _14839_ (.B1(_08323_),
    .Y(_01510_),
    .A1(net279),
    .A2(net496));
 sg13g2_buf_1 fanout176 (.A(_07719_),
    .X(net176));
 sg13g2_nand2_1 _14841_ (.Y(_08325_),
    .A(\dp.rf.rf[7][9] ),
    .B(net495));
 sg13g2_o21ai_1 _14842_ (.B1(_08325_),
    .Y(_01511_),
    .A1(net275),
    .A2(net495));
 sg13g2_nand2_1 _14843_ (.Y(_08326_),
    .A(\dp.rf.rf[7][10] ),
    .B(net494));
 sg13g2_o21ai_1 _14844_ (.B1(_08326_),
    .Y(_01512_),
    .A1(net266),
    .A2(net494));
 sg13g2_buf_1 fanout175 (.A(net176),
    .X(net175));
 sg13g2_nand2_1 _14846_ (.Y(_08328_),
    .A(\dp.rf.rf[7][11] ),
    .B(net497));
 sg13g2_o21ai_1 _14847_ (.B1(_08328_),
    .Y(_01513_),
    .A1(net263),
    .A2(net496));
 sg13g2_nand2_1 _14848_ (.Y(_08329_),
    .A(\dp.rf.rf[7][12] ),
    .B(net494));
 sg13g2_o21ai_1 _14849_ (.B1(_08329_),
    .Y(_01514_),
    .A1(net259),
    .A2(net494));
 sg13g2_mux2_1 _14850_ (.A0(net252),
    .A1(\dp.rf.rf[7][13] ),
    .S(net495),
    .X(_01515_));
 sg13g2_nand2_1 _14851_ (.Y(_08330_),
    .A(\dp.rf.rf[7][14] ),
    .B(net490));
 sg13g2_o21ai_1 _14852_ (.B1(_08330_),
    .Y(_01516_),
    .A1(net245),
    .A2(net490));
 sg13g2_nand2_1 _14853_ (.Y(_08331_),
    .A(\dp.rf.rf[7][15] ),
    .B(net493));
 sg13g2_o21ai_1 _14854_ (.B1(_08331_),
    .Y(_01517_),
    .A1(net243),
    .A2(net493));
 sg13g2_nand2_1 _14855_ (.Y(_08332_),
    .A(\dp.rf.rf[7][16] ),
    .B(net493));
 sg13g2_o21ai_1 _14856_ (.B1(_08332_),
    .Y(_01518_),
    .A1(net238),
    .A2(net493));
 sg13g2_nand2_1 _14857_ (.Y(_08333_),
    .A(\dp.rf.rf[7][17] ),
    .B(net492));
 sg13g2_o21ai_1 _14858_ (.B1(_08333_),
    .Y(_01519_),
    .A1(net232),
    .A2(net492));
 sg13g2_nand2_1 _14859_ (.Y(_08334_),
    .A(\dp.rf.rf[7][18] ),
    .B(net495));
 sg13g2_o21ai_1 _14860_ (.B1(_08334_),
    .Y(_01520_),
    .A1(net227),
    .A2(net495));
 sg13g2_nand2_1 _14861_ (.Y(_08335_),
    .A(\dp.rf.rf[7][19] ),
    .B(net488));
 sg13g2_o21ai_1 _14862_ (.B1(_08335_),
    .Y(_01521_),
    .A1(net223),
    .A2(net488));
 sg13g2_buf_2 fanout174 (.A(net175),
    .X(net174));
 sg13g2_nand2_1 _14864_ (.Y(_08337_),
    .A(\dp.rf.rf[7][20] ),
    .B(net491));
 sg13g2_o21ai_1 _14865_ (.B1(_08337_),
    .Y(_01522_),
    .A1(net214),
    .A2(net491));
 sg13g2_nand2_1 _14866_ (.Y(_08338_),
    .A(\dp.rf.rf[7][21] ),
    .B(net489));
 sg13g2_o21ai_1 _14867_ (.B1(_08338_),
    .Y(_01523_),
    .A1(net209),
    .A2(net489));
 sg13g2_buf_2 fanout173 (.A(_07731_),
    .X(net173));
 sg13g2_nand2_1 _14869_ (.Y(_08340_),
    .A(\dp.rf.rf[7][22] ),
    .B(net491));
 sg13g2_o21ai_1 _14870_ (.B1(_08340_),
    .Y(_01524_),
    .A1(net206),
    .A2(net491));
 sg13g2_nand2_1 _14871_ (.Y(_08341_),
    .A(\dp.rf.rf[7][23] ),
    .B(net488));
 sg13g2_o21ai_1 _14872_ (.B1(_08341_),
    .Y(_01525_),
    .A1(net202),
    .A2(net488));
 sg13g2_nand2_1 _14873_ (.Y(_08342_),
    .A(\dp.rf.rf[7][24] ),
    .B(net489));
 sg13g2_o21ai_1 _14874_ (.B1(_08342_),
    .Y(_01526_),
    .A1(net196),
    .A2(net489));
 sg13g2_nand2_1 _14875_ (.Y(_08343_),
    .A(\dp.rf.rf[7][25] ),
    .B(net489));
 sg13g2_o21ai_1 _14876_ (.B1(_08343_),
    .Y(_01527_),
    .A1(net191),
    .A2(net489));
 sg13g2_nand2_1 _14877_ (.Y(_08344_),
    .A(\dp.rf.rf[7][26] ),
    .B(net491));
 sg13g2_o21ai_1 _14878_ (.B1(_08344_),
    .Y(_01528_),
    .A1(net187),
    .A2(net491));
 sg13g2_nand2_1 _14879_ (.Y(_08345_),
    .A(\dp.rf.rf[7][27] ),
    .B(net488));
 sg13g2_o21ai_1 _14880_ (.B1(_08345_),
    .Y(_01529_),
    .A1(net182),
    .A2(net488));
 sg13g2_nand2_1 _14881_ (.Y(_08346_),
    .A(\dp.rf.rf[7][28] ),
    .B(net489));
 sg13g2_o21ai_1 _14882_ (.B1(_08346_),
    .Y(_01530_),
    .A1(net305),
    .A2(net489));
 sg13g2_nand2_1 _14883_ (.Y(_08347_),
    .A(\dp.rf.rf[7][29] ),
    .B(net492));
 sg13g2_o21ai_1 _14884_ (.B1(_08347_),
    .Y(_01531_),
    .A1(net178),
    .A2(net492));
 sg13g2_nand2_1 _14885_ (.Y(_08348_),
    .A(\dp.rf.rf[7][30] ),
    .B(net491));
 sg13g2_o21ai_1 _14886_ (.B1(_08348_),
    .Y(_01532_),
    .A1(net170),
    .A2(net491));
 sg13g2_nand2_1 _14887_ (.Y(_08349_),
    .A(\dp.rf.rf[7][31] ),
    .B(net488));
 sg13g2_o21ai_1 _14888_ (.B1(_08349_),
    .Y(_01533_),
    .A1(net168),
    .A2(net488));
 sg13g2_buf_2 fanout172 (.A(_07731_),
    .X(net172));
 sg13g2_buf_2 fanout171 (.A(_07731_),
    .X(net171));
 sg13g2_buf_2 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_1 fanout169 (.A(_07741_),
    .X(net169));
 sg13g2_buf_2 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_2 fanout167 (.A(net169),
    .X(net167));
 sg13g2_buf_2 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_2 fanout165 (.A(net167),
    .X(net165));
 sg13g2_buf_1 output164 (.A(net164),
    .X(writedata[9]));
 sg13g2_buf_1 output163 (.A(net163),
    .X(writedata[8]));
 sg13g2_buf_1 output162 (.A(net162),
    .X(writedata[7]));
 sg13g2_buf_1 output161 (.A(net161),
    .X(writedata[6]));
 sg13g2_buf_1 output160 (.A(net160),
    .X(writedata[5]));
 sg13g2_buf_1 output159 (.A(net159),
    .X(writedata[4]));
 sg13g2_buf_1 output158 (.A(net158),
    .X(writedata[3]));
 sg13g2_buf_1 output157 (.A(net157),
    .X(writedata[31]));
 sg13g2_buf_1 output156 (.A(net156),
    .X(writedata[30]));
 sg13g2_buf_1 output155 (.A(net155),
    .X(writedata[2]));
 sg13g2_buf_1 output154 (.A(net154),
    .X(writedata[29]));
 sg13g2_buf_1 output153 (.A(net153),
    .X(writedata[28]));
 sg13g2_buf_1 output152 (.A(net152),
    .X(writedata[27]));
 sg13g2_buf_1 output151 (.A(net151),
    .X(writedata[26]));
 sg13g2_buf_1 output150 (.A(net150),
    .X(writedata[25]));
 sg13g2_buf_1 output149 (.A(net149),
    .X(writedata[24]));
 sg13g2_buf_1 output148 (.A(net148),
    .X(writedata[23]));
 sg13g2_buf_1 output147 (.A(net147),
    .X(writedata[22]));
 sg13g2_buf_1 output146 (.A(net146),
    .X(writedata[21]));
 sg13g2_buf_1 output145 (.A(net145),
    .X(writedata[20]));
 sg13g2_buf_1 output144 (.A(net144),
    .X(writedata[1]));
 sg13g2_buf_1 output143 (.A(net143),
    .X(writedata[19]));
 sg13g2_nand2_1 _14919_ (.Y(_08350_),
    .A(_07841_),
    .B(_08311_));
 sg13g2_buf_1 output142 (.A(net142),
    .X(writedata[18]));
 sg13g2_buf_1 output141 (.A(net141),
    .X(writedata[17]));
 sg13g2_buf_1 output140 (.A(net140),
    .X(writedata[16]));
 sg13g2_nand2_1 _14923_ (.Y(_08354_),
    .A(\dp.rf.rf[4][0] ),
    .B(net725));
 sg13g2_o21ai_1 _14924_ (.B1(_08354_),
    .Y(_01564_),
    .A1(net303),
    .A2(net725));
 sg13g2_nand2_1 _14925_ (.Y(_08355_),
    .A(\dp.rf.rf[4][1] ),
    .B(net726));
 sg13g2_o21ai_1 _14926_ (.B1(_08355_),
    .Y(_01565_),
    .A1(net297),
    .A2(net726));
 sg13g2_nand2_1 _14927_ (.Y(_08356_),
    .A(\dp.rf.rf[4][2] ),
    .B(net726));
 sg13g2_o21ai_1 _14928_ (.B1(_08356_),
    .Y(_01566_),
    .A1(net320),
    .A2(net726));
 sg13g2_nand2_1 _14929_ (.Y(_08357_),
    .A(\dp.rf.rf[4][3] ),
    .B(net727));
 sg13g2_o21ai_1 _14930_ (.B1(_08357_),
    .Y(_01567_),
    .A1(net316),
    .A2(net726));
 sg13g2_mux2_1 _14931_ (.A0(net291),
    .A1(\dp.rf.rf[4][4] ),
    .S(net725),
    .X(_01568_));
 sg13g2_nand2_1 _14932_ (.Y(_08358_),
    .A(\dp.rf.rf[4][5] ),
    .B(net724));
 sg13g2_o21ai_1 _14933_ (.B1(_08358_),
    .Y(_01569_),
    .A1(net311),
    .A2(net723));
 sg13g2_nand2_1 _14934_ (.Y(_08359_),
    .A(\dp.rf.rf[4][6] ),
    .B(net723));
 sg13g2_o21ai_1 _14935_ (.B1(_08359_),
    .Y(_01570_),
    .A1(net285),
    .A2(net723));
 sg13g2_nand2_1 _14936_ (.Y(_08360_),
    .A(\dp.rf.rf[4][7] ),
    .B(net724));
 sg13g2_o21ai_1 _14937_ (.B1(_08360_),
    .Y(_01571_),
    .A1(net283),
    .A2(net723));
 sg13g2_nand2_1 _14938_ (.Y(_08361_),
    .A(\dp.rf.rf[4][8] ),
    .B(net726));
 sg13g2_o21ai_1 _14939_ (.B1(_08361_),
    .Y(_01572_),
    .A1(net279),
    .A2(net726));
 sg13g2_buf_1 output139 (.A(net139),
    .X(writedata[15]));
 sg13g2_nand2_1 _14941_ (.Y(_08363_),
    .A(\dp.rf.rf[4][9] ),
    .B(net725));
 sg13g2_o21ai_1 _14942_ (.B1(_08363_),
    .Y(_01573_),
    .A1(net275),
    .A2(net725));
 sg13g2_nand2_1 _14943_ (.Y(_08364_),
    .A(\dp.rf.rf[4][10] ),
    .B(net724));
 sg13g2_o21ai_1 _14944_ (.B1(_08364_),
    .Y(_01574_),
    .A1(net267),
    .A2(net724));
 sg13g2_buf_1 output138 (.A(net138),
    .X(writedata[14]));
 sg13g2_nand2_1 _14946_ (.Y(_08366_),
    .A(\dp.rf.rf[4][11] ),
    .B(net726));
 sg13g2_o21ai_1 _14947_ (.B1(_08366_),
    .Y(_01575_),
    .A1(net263),
    .A2(net727));
 sg13g2_nand2_1 _14948_ (.Y(_08367_),
    .A(\dp.rf.rf[4][12] ),
    .B(net724));
 sg13g2_o21ai_1 _14949_ (.B1(_08367_),
    .Y(_01576_),
    .A1(net259),
    .A2(net724));
 sg13g2_mux2_1 _14950_ (.A0(net250),
    .A1(\dp.rf.rf[4][13] ),
    .S(net725),
    .X(_01577_));
 sg13g2_nand2_1 _14951_ (.Y(_08368_),
    .A(\dp.rf.rf[4][14] ),
    .B(net718));
 sg13g2_o21ai_1 _14952_ (.B1(_08368_),
    .Y(_01578_),
    .A1(net245),
    .A2(net718));
 sg13g2_nand2_1 _14953_ (.Y(_08369_),
    .A(\dp.rf.rf[4][15] ),
    .B(net723));
 sg13g2_o21ai_1 _14954_ (.B1(_08369_),
    .Y(_01579_),
    .A1(net243),
    .A2(net723));
 sg13g2_nand2_1 _14955_ (.Y(_08370_),
    .A(\dp.rf.rf[4][16] ),
    .B(net723));
 sg13g2_o21ai_1 _14956_ (.B1(_08370_),
    .Y(_01580_),
    .A1(net236),
    .A2(net723));
 sg13g2_nand2_1 _14957_ (.Y(_08371_),
    .A(\dp.rf.rf[4][17] ),
    .B(net721));
 sg13g2_o21ai_1 _14958_ (.B1(_08371_),
    .Y(_01581_),
    .A1(net230),
    .A2(net721));
 sg13g2_nand2_1 _14959_ (.Y(_08372_),
    .A(\dp.rf.rf[4][18] ),
    .B(net725));
 sg13g2_o21ai_1 _14960_ (.B1(_08372_),
    .Y(_01582_),
    .A1(net225),
    .A2(net725));
 sg13g2_nand2_1 _14961_ (.Y(_08373_),
    .A(\dp.rf.rf[4][19] ),
    .B(net722));
 sg13g2_o21ai_1 _14962_ (.B1(_08373_),
    .Y(_01583_),
    .A1(net223),
    .A2(net722));
 sg13g2_buf_1 output137 (.A(net137),
    .X(writedata[13]));
 sg13g2_nand2_1 _14964_ (.Y(_08375_),
    .A(\dp.rf.rf[4][20] ),
    .B(net720));
 sg13g2_o21ai_1 _14965_ (.B1(_08375_),
    .Y(_01584_),
    .A1(net214),
    .A2(net720));
 sg13g2_nand2_1 _14966_ (.Y(_08376_),
    .A(\dp.rf.rf[4][21] ),
    .B(net719));
 sg13g2_o21ai_1 _14967_ (.B1(_08376_),
    .Y(_01585_),
    .A1(net210),
    .A2(net719));
 sg13g2_buf_1 output136 (.A(net136),
    .X(writedata[12]));
 sg13g2_nand2_1 _14969_ (.Y(_08378_),
    .A(\dp.rf.rf[4][22] ),
    .B(net720));
 sg13g2_o21ai_1 _14970_ (.B1(_08378_),
    .Y(_01586_),
    .A1(net205),
    .A2(net720));
 sg13g2_nand2_1 _14971_ (.Y(_08379_),
    .A(\dp.rf.rf[4][23] ),
    .B(net718));
 sg13g2_o21ai_1 _14972_ (.B1(_08379_),
    .Y(_01587_),
    .A1(net202),
    .A2(net718));
 sg13g2_nand2_1 _14973_ (.Y(_08380_),
    .A(\dp.rf.rf[4][24] ),
    .B(net719));
 sg13g2_o21ai_1 _14974_ (.B1(_08380_),
    .Y(_01588_),
    .A1(net195),
    .A2(net719));
 sg13g2_nand2_1 _14975_ (.Y(_08381_),
    .A(\dp.rf.rf[4][25] ),
    .B(net719));
 sg13g2_o21ai_1 _14976_ (.B1(_08381_),
    .Y(_01589_),
    .A1(net191),
    .A2(net719));
 sg13g2_nand2_1 _14977_ (.Y(_08382_),
    .A(\dp.rf.rf[4][26] ),
    .B(net720));
 sg13g2_o21ai_1 _14978_ (.B1(_08382_),
    .Y(_01590_),
    .A1(net186),
    .A2(net720));
 sg13g2_nand2_1 _14979_ (.Y(_08383_),
    .A(\dp.rf.rf[4][27] ),
    .B(net718));
 sg13g2_o21ai_1 _14980_ (.B1(_08383_),
    .Y(_01591_),
    .A1(net182),
    .A2(net718));
 sg13g2_nand2_1 _14981_ (.Y(_08384_),
    .A(\dp.rf.rf[4][28] ),
    .B(net719));
 sg13g2_o21ai_1 _14982_ (.B1(_08384_),
    .Y(_01592_),
    .A1(net305),
    .A2(net719));
 sg13g2_nand2_1 _14983_ (.Y(_08385_),
    .A(\dp.rf.rf[4][29] ),
    .B(net721));
 sg13g2_o21ai_1 _14984_ (.B1(_08385_),
    .Y(_01593_),
    .A1(net178),
    .A2(net721));
 sg13g2_nand2_1 _14985_ (.Y(_08386_),
    .A(\dp.rf.rf[4][30] ),
    .B(net720));
 sg13g2_o21ai_1 _14986_ (.B1(_08386_),
    .Y(_01594_),
    .A1(net170),
    .A2(net720));
 sg13g2_nand2_1 _14987_ (.Y(_08387_),
    .A(\dp.rf.rf[4][31] ),
    .B(net718));
 sg13g2_o21ai_1 _14988_ (.B1(_08387_),
    .Y(_01595_),
    .A1(net167),
    .A2(net718));
 sg13g2_buf_1 output135 (.A(net135),
    .X(writedata[11]));
 sg13g2_nand2_1 _14990_ (.Y(_08389_),
    .A(_07746_),
    .B(_07795_));
 sg13g2_buf_1 output134 (.A(net134),
    .X(writedata[10]));
 sg13g2_buf_1 output133 (.A(net133),
    .X(writedata[0]));
 sg13g2_buf_1 output132 (.A(net132),
    .X(suspend));
 sg13g2_nand2_1 _14994_ (.Y(_08393_),
    .A(\dp.rf.rf[9][0] ),
    .B(net485));
 sg13g2_o21ai_1 _14995_ (.B1(_08393_),
    .Y(_01596_),
    .A1(net300),
    .A2(net485));
 sg13g2_nand2_1 _14996_ (.Y(_08394_),
    .A(\dp.rf.rf[9][1] ),
    .B(net487));
 sg13g2_o21ai_1 _14997_ (.B1(_08394_),
    .Y(_01597_),
    .A1(net295),
    .A2(net487));
 sg13g2_nand2_1 _14998_ (.Y(_08395_),
    .A(\dp.rf.rf[9][2] ),
    .B(net487));
 sg13g2_o21ai_1 _14999_ (.B1(_08395_),
    .Y(_01598_),
    .A1(net320),
    .A2(net486));
 sg13g2_nand2_1 _15000_ (.Y(_08396_),
    .A(\dp.rf.rf[9][3] ),
    .B(net486));
 sg13g2_o21ai_1 _15001_ (.B1(_08396_),
    .Y(_01599_),
    .A1(net317),
    .A2(net486));
 sg13g2_mux2_1 _15002_ (.A0(net294),
    .A1(\dp.rf.rf[9][4] ),
    .S(net485),
    .X(_01600_));
 sg13g2_nand2_1 _15003_ (.Y(_08397_),
    .A(\dp.rf.rf[9][5] ),
    .B(net483));
 sg13g2_o21ai_1 _15004_ (.B1(_08397_),
    .Y(_01601_),
    .A1(net310),
    .A2(net483));
 sg13g2_nand2_1 _15005_ (.Y(_08398_),
    .A(\dp.rf.rf[9][6] ),
    .B(net483));
 sg13g2_o21ai_1 _15006_ (.B1(_08398_),
    .Y(_01602_),
    .A1(net286),
    .A2(net483));
 sg13g2_nand2_1 _15007_ (.Y(_08399_),
    .A(\dp.rf.rf[9][7] ),
    .B(net483));
 sg13g2_o21ai_1 _15008_ (.B1(_08399_),
    .Y(_01603_),
    .A1(net281),
    .A2(net483));
 sg13g2_nand2_1 _15009_ (.Y(_08400_),
    .A(\dp.rf.rf[9][8] ),
    .B(net486));
 sg13g2_o21ai_1 _15010_ (.B1(_08400_),
    .Y(_01604_),
    .A1(net276),
    .A2(net484));
 sg13g2_buf_1 output131 (.A(net131),
    .X(pc[9]));
 sg13g2_nand2_1 _15012_ (.Y(_08402_),
    .A(\dp.rf.rf[9][9] ),
    .B(net485));
 sg13g2_o21ai_1 _15013_ (.B1(_08402_),
    .Y(_01605_),
    .A1(net274),
    .A2(net485));
 sg13g2_nand2_1 _15014_ (.Y(_08403_),
    .A(\dp.rf.rf[9][10] ),
    .B(net484));
 sg13g2_o21ai_1 _15015_ (.B1(_08403_),
    .Y(_01606_),
    .A1(net266),
    .A2(net484));
 sg13g2_buf_1 output130 (.A(net130),
    .X(pc[8]));
 sg13g2_nand2_1 _15017_ (.Y(_08405_),
    .A(\dp.rf.rf[9][11] ),
    .B(net486));
 sg13g2_o21ai_1 _15018_ (.B1(_08405_),
    .Y(_01607_),
    .A1(net260),
    .A2(net486));
 sg13g2_nand2_1 _15019_ (.Y(_08406_),
    .A(\dp.rf.rf[9][12] ),
    .B(net484));
 sg13g2_o21ai_1 _15020_ (.B1(_08406_),
    .Y(_01608_),
    .A1(net254),
    .A2(net484));
 sg13g2_mux2_1 _15021_ (.A0(net249),
    .A1(\dp.rf.rf[9][13] ),
    .S(net485),
    .X(_01609_));
 sg13g2_nand2_1 _15022_ (.Y(_08407_),
    .A(\dp.rf.rf[9][14] ),
    .B(net480));
 sg13g2_o21ai_1 _15023_ (.B1(_08407_),
    .Y(_01610_),
    .A1(net247),
    .A2(net479));
 sg13g2_nand2_1 _15024_ (.Y(_08408_),
    .A(\dp.rf.rf[9][15] ),
    .B(net483));
 sg13g2_o21ai_1 _15025_ (.B1(_08408_),
    .Y(_01611_),
    .A1(net244),
    .A2(net483));
 sg13g2_nand2_1 _15026_ (.Y(_08409_),
    .A(\dp.rf.rf[9][16] ),
    .B(net484));
 sg13g2_o21ai_1 _15027_ (.B1(_08409_),
    .Y(_01612_),
    .A1(net238),
    .A2(net484));
 sg13g2_buf_1 output129 (.A(net129),
    .X(pc[7]));
 sg13g2_nand2_1 _15029_ (.Y(_08411_),
    .A(\dp.rf.rf[9][17] ),
    .B(net479));
 sg13g2_o21ai_1 _15030_ (.B1(_08411_),
    .Y(_01613_),
    .A1(net229),
    .A2(net480));
 sg13g2_nand2_1 _15031_ (.Y(_08412_),
    .A(\dp.rf.rf[9][18] ),
    .B(net485));
 sg13g2_o21ai_1 _15032_ (.B1(_08412_),
    .Y(_01614_),
    .A1(net227),
    .A2(net485));
 sg13g2_nand2_1 _15033_ (.Y(_08413_),
    .A(\dp.rf.rf[9][19] ),
    .B(net479));
 sg13g2_o21ai_1 _15034_ (.B1(_08413_),
    .Y(_01615_),
    .A1(net220),
    .A2(net479));
 sg13g2_buf_1 output128 (.A(net128),
    .X(pc[6]));
 sg13g2_nand2_1 _15036_ (.Y(_08415_),
    .A(\dp.rf.rf[9][20] ),
    .B(net481));
 sg13g2_o21ai_1 _15037_ (.B1(_08415_),
    .Y(_01616_),
    .A1(net214),
    .A2(net481));
 sg13g2_nand2_1 _15038_ (.Y(_08416_),
    .A(\dp.rf.rf[9][21] ),
    .B(net480));
 sg13g2_o21ai_1 _15039_ (.B1(_08416_),
    .Y(_01617_),
    .A1(net209),
    .A2(net478));
 sg13g2_buf_1 output127 (.A(net127),
    .X(pc[5]));
 sg13g2_nand2_1 _15041_ (.Y(_08418_),
    .A(\dp.rf.rf[9][22] ),
    .B(net482));
 sg13g2_o21ai_1 _15042_ (.B1(_08418_),
    .Y(_01618_),
    .A1(net206),
    .A2(net482));
 sg13g2_nand2_1 _15043_ (.Y(_08419_),
    .A(\dp.rf.rf[9][23] ),
    .B(net479));
 sg13g2_o21ai_1 _15044_ (.B1(_08419_),
    .Y(_01619_),
    .A1(net203),
    .A2(net479));
 sg13g2_nand2_1 _15045_ (.Y(_08420_),
    .A(\dp.rf.rf[9][24] ),
    .B(net478));
 sg13g2_o21ai_1 _15046_ (.B1(_08420_),
    .Y(_01620_),
    .A1(net199),
    .A2(net478));
 sg13g2_nand2_1 _15047_ (.Y(_08421_),
    .A(\dp.rf.rf[9][25] ),
    .B(net478));
 sg13g2_o21ai_1 _15048_ (.B1(_08421_),
    .Y(_01621_),
    .A1(net192),
    .A2(net478));
 sg13g2_nand2_1 _15049_ (.Y(_08422_),
    .A(\dp.rf.rf[9][26] ),
    .B(net481));
 sg13g2_o21ai_1 _15050_ (.B1(_08422_),
    .Y(_01622_),
    .A1(net187),
    .A2(net481));
 sg13g2_nand2_1 _15051_ (.Y(_08423_),
    .A(\dp.rf.rf[9][27] ),
    .B(net478));
 sg13g2_o21ai_1 _15052_ (.B1(_08423_),
    .Y(_01623_),
    .A1(net181),
    .A2(net478));
 sg13g2_nand2_1 _15053_ (.Y(_08424_),
    .A(\dp.rf.rf[9][28] ),
    .B(net478));
 sg13g2_o21ai_1 _15054_ (.B1(_08424_),
    .Y(_01624_),
    .A1(net307),
    .A2(net480));
 sg13g2_nand2_1 _15055_ (.Y(_08425_),
    .A(\dp.rf.rf[9][29] ),
    .B(net481));
 sg13g2_o21ai_1 _15056_ (.B1(_08425_),
    .Y(_01625_),
    .A1(net177),
    .A2(net481));
 sg13g2_buf_1 output126 (.A(net126),
    .X(pc[4]));
 sg13g2_nand2_1 _15058_ (.Y(_08427_),
    .A(\dp.rf.rf[9][30] ),
    .B(net481));
 sg13g2_o21ai_1 _15059_ (.B1(_08427_),
    .Y(_01626_),
    .A1(net170),
    .A2(net481));
 sg13g2_nand2_1 _15060_ (.Y(_08428_),
    .A(\dp.rf.rf[9][31] ),
    .B(net479));
 sg13g2_o21ai_1 _15061_ (.B1(_08428_),
    .Y(_01627_),
    .A1(net168),
    .A2(net479));
 sg13g2_nand2_1 _15062_ (.Y(_08429_),
    .A(_07930_),
    .B(_08191_));
 sg13g2_buf_1 output125 (.A(net125),
    .X(pc[3]));
 sg13g2_buf_1 output124 (.A(net124),
    .X(pc[31]));
 sg13g2_buf_1 output123 (.A(net123),
    .X(pc[30]));
 sg13g2_nand2_1 _15066_ (.Y(_08433_),
    .A(\dp.rf.rf[22][0] ),
    .B(net711));
 sg13g2_o21ai_1 _15067_ (.B1(_08433_),
    .Y(_01628_),
    .A1(net301),
    .A2(net711));
 sg13g2_nand2_1 _15068_ (.Y(_08434_),
    .A(\dp.rf.rf[22][1] ),
    .B(net715));
 sg13g2_o21ai_1 _15069_ (.B1(_08434_),
    .Y(_01629_),
    .A1(net297),
    .A2(net715));
 sg13g2_buf_1 output122 (.A(net122),
    .X(pc[2]));
 sg13g2_nand2_1 _15071_ (.Y(_08436_),
    .A(\dp.rf.rf[22][2] ),
    .B(net716));
 sg13g2_o21ai_1 _15072_ (.B1(_08436_),
    .Y(_01630_),
    .A1(net324),
    .A2(net715));
 sg13g2_nand2_1 _15073_ (.Y(_08437_),
    .A(\dp.rf.rf[22][3] ),
    .B(net715));
 sg13g2_o21ai_1 _15074_ (.B1(_08437_),
    .Y(_01631_),
    .A1(net319),
    .A2(net715));
 sg13g2_nor2_2 _15075_ (.A(_07924_),
    .B(_08201_),
    .Y(_08438_));
 sg13g2_buf_1 output121 (.A(net121),
    .X(pc[29]));
 sg13g2_mux2_1 _15077_ (.A0(\dp.rf.rf[22][4] ),
    .A1(net293),
    .S(_08438_),
    .X(_01632_));
 sg13g2_nand2_1 _15078_ (.Y(_08440_),
    .A(\dp.rf.rf[22][5] ),
    .B(net714));
 sg13g2_o21ai_1 _15079_ (.B1(_08440_),
    .Y(_01633_),
    .A1(net313),
    .A2(net714));
 sg13g2_nand2_1 _15080_ (.Y(_08441_),
    .A(\dp.rf.rf[22][6] ),
    .B(net714));
 sg13g2_o21ai_1 _15081_ (.B1(_08441_),
    .Y(_01634_),
    .A1(net287),
    .A2(net714));
 sg13g2_nand2_1 _15082_ (.Y(_08442_),
    .A(\dp.rf.rf[22][7] ),
    .B(net713));
 sg13g2_o21ai_1 _15083_ (.B1(_08442_),
    .Y(_01635_),
    .A1(net281),
    .A2(net713));
 sg13g2_nand2_1 _15084_ (.Y(_08443_),
    .A(\dp.rf.rf[22][8] ),
    .B(net716));
 sg13g2_o21ai_1 _15085_ (.B1(_08443_),
    .Y(_01636_),
    .A1(net277),
    .A2(net716));
 sg13g2_nand2_1 _15086_ (.Y(_08444_),
    .A(\dp.rf.rf[22][9] ),
    .B(net713));
 sg13g2_o21ai_1 _15087_ (.B1(_08444_),
    .Y(_01637_),
    .A1(net271),
    .A2(net713));
 sg13g2_nand2_1 _15088_ (.Y(_08445_),
    .A(\dp.rf.rf[22][10] ),
    .B(net715));
 sg13g2_o21ai_1 _15089_ (.B1(_08445_),
    .Y(_01638_),
    .A1(net268),
    .A2(net715));
 sg13g2_buf_1 output120 (.A(net120),
    .X(pc[28]));
 sg13g2_nand2_1 _15091_ (.Y(_08447_),
    .A(\dp.rf.rf[22][11] ),
    .B(net715));
 sg13g2_o21ai_1 _15092_ (.B1(_08447_),
    .Y(_01639_),
    .A1(net264),
    .A2(net716));
 sg13g2_nand2_1 _15093_ (.Y(_08448_),
    .A(\dp.rf.rf[22][12] ),
    .B(net714));
 sg13g2_o21ai_1 _15094_ (.B1(_08448_),
    .Y(_01640_),
    .A1(net257),
    .A2(net714));
 sg13g2_mux2_1 _15095_ (.A0(\dp.rf.rf[22][13] ),
    .A1(net252),
    .S(_08438_),
    .X(_01641_));
 sg13g2_buf_1 output119 (.A(net119),
    .X(pc[27]));
 sg13g2_nand2_1 _15097_ (.Y(_08450_),
    .A(\dp.rf.rf[22][14] ),
    .B(net710));
 sg13g2_o21ai_1 _15098_ (.B1(_08450_),
    .Y(_01642_),
    .A1(net245),
    .A2(net710));
 sg13g2_nand2_1 _15099_ (.Y(_08451_),
    .A(\dp.rf.rf[22][15] ),
    .B(net713));
 sg13g2_o21ai_1 _15100_ (.B1(_08451_),
    .Y(_01643_),
    .A1(net240),
    .A2(net713));
 sg13g2_nand2_1 _15101_ (.Y(_08452_),
    .A(\dp.rf.rf[22][16] ),
    .B(net713));
 sg13g2_o21ai_1 _15102_ (.B1(_08452_),
    .Y(_01644_),
    .A1(net237),
    .A2(net713));
 sg13g2_nand2_1 _15103_ (.Y(_08453_),
    .A(\dp.rf.rf[22][17] ),
    .B(net717));
 sg13g2_o21ai_1 _15104_ (.B1(_08453_),
    .Y(_01645_),
    .A1(net232),
    .A2(net712));
 sg13g2_nand2_1 _15105_ (.Y(_08454_),
    .A(\dp.rf.rf[22][18] ),
    .B(net711));
 sg13g2_o21ai_1 _15106_ (.B1(_08454_),
    .Y(_01646_),
    .A1(net224),
    .A2(net711));
 sg13g2_nand2_1 _15107_ (.Y(_08455_),
    .A(\dp.rf.rf[22][19] ),
    .B(net712));
 sg13g2_o21ai_1 _15108_ (.B1(_08455_),
    .Y(_01647_),
    .A1(net221),
    .A2(net712));
 sg13g2_nand2_1 _15109_ (.Y(_08456_),
    .A(\dp.rf.rf[22][20] ),
    .B(net710));
 sg13g2_o21ai_1 _15110_ (.B1(_08456_),
    .Y(_01648_),
    .A1(net216),
    .A2(net710));
 sg13g2_nand2_1 _15111_ (.Y(_08457_),
    .A(\dp.rf.rf[22][21] ),
    .B(net710));
 sg13g2_o21ai_1 _15112_ (.B1(_08457_),
    .Y(_01649_),
    .A1(net211),
    .A2(net710));
 sg13g2_nor2_1 _15113_ (.A(\dp.rf.rf[22][22] ),
    .B(_08438_),
    .Y(_08458_));
 sg13g2_a21oi_1 _15114_ (.A1(net208),
    .A2(_08438_),
    .Y(_01650_),
    .B1(_08458_));
 sg13g2_nand2_1 _15115_ (.Y(_08459_),
    .A(\dp.rf.rf[22][23] ),
    .B(net709));
 sg13g2_o21ai_1 _15116_ (.B1(_08459_),
    .Y(_01651_),
    .A1(net200),
    .A2(net709));
 sg13g2_nand2_1 _15117_ (.Y(_08460_),
    .A(\dp.rf.rf[22][24] ),
    .B(net712));
 sg13g2_o21ai_1 _15118_ (.B1(_08460_),
    .Y(_01652_),
    .A1(net198),
    .A2(net712));
 sg13g2_nand2_1 _15119_ (.Y(_08461_),
    .A(\dp.rf.rf[22][25] ),
    .B(net709));
 sg13g2_o21ai_1 _15120_ (.B1(_08461_),
    .Y(_01653_),
    .A1(net189),
    .A2(net709));
 sg13g2_nand2_1 _15121_ (.Y(_08462_),
    .A(\dp.rf.rf[22][26] ),
    .B(net709));
 sg13g2_o21ai_1 _15122_ (.B1(_08462_),
    .Y(_01654_),
    .A1(net183),
    .A2(net709));
 sg13g2_nand2_1 _15123_ (.Y(_08463_),
    .A(\dp.rf.rf[22][27] ),
    .B(net709));
 sg13g2_o21ai_1 _15124_ (.B1(_08463_),
    .Y(_01655_),
    .A1(net179),
    .A2(net709));
 sg13g2_nand2_1 _15125_ (.Y(_08464_),
    .A(\dp.rf.rf[22][28] ),
    .B(net710));
 sg13g2_o21ai_1 _15126_ (.B1(_08464_),
    .Y(_01656_),
    .A1(net306),
    .A2(net710));
 sg13g2_nor2_1 _15127_ (.A(\dp.rf.rf[22][29] ),
    .B(_08438_),
    .Y(_08465_));
 sg13g2_a21oi_1 _15128_ (.A1(net174),
    .A2(_08438_),
    .Y(_01657_),
    .B1(_08465_));
 sg13g2_nand2_1 _15129_ (.Y(_08466_),
    .A(\dp.rf.rf[22][30] ),
    .B(net712));
 sg13g2_o21ai_1 _15130_ (.B1(_08466_),
    .Y(_01658_),
    .A1(net172),
    .A2(net712));
 sg13g2_nand2_1 _15131_ (.Y(_08467_),
    .A(\dp.rf.rf[22][31] ),
    .B(net711));
 sg13g2_o21ai_1 _15132_ (.B1(_08467_),
    .Y(_01659_),
    .A1(net165),
    .A2(net711));
 sg13g2_nand2_2 _15133_ (.Y(_08468_),
    .A(net1247),
    .B(_07745_));
 sg13g2_buf_1 output118 (.A(net118),
    .X(pc[26]));
 sg13g2_nor2_1 _15135_ (.A(_07790_),
    .B(_08468_),
    .Y(_08470_));
 sg13g2_buf_1 output117 (.A(net117),
    .X(pc[25]));
 sg13g2_buf_1 output116 (.A(net116),
    .X(pc[24]));
 sg13g2_nor2_1 _15138_ (.A(\dp.rf.rf[25][0] ),
    .B(_08470_),
    .Y(_08473_));
 sg13g2_a21oi_1 _15139_ (.A1(net302),
    .A2(net477),
    .Y(_01660_),
    .B1(_08473_));
 sg13g2_or2_1 _15140_ (.X(_08474_),
    .B(_08468_),
    .A(_07790_));
 sg13g2_buf_1 output115 (.A(net115),
    .X(pc[23]));
 sg13g2_buf_1 output114 (.A(net114),
    .X(pc[22]));
 sg13g2_buf_1 output113 (.A(net113),
    .X(pc[21]));
 sg13g2_nand2_1 _15144_ (.Y(_08478_),
    .A(\dp.rf.rf[25][1] ),
    .B(net474));
 sg13g2_o21ai_1 _15145_ (.B1(_08478_),
    .Y(_01661_),
    .A1(net298),
    .A2(net473));
 sg13g2_nand2_1 _15146_ (.Y(_08479_),
    .A(\dp.rf.rf[25][2] ),
    .B(net473));
 sg13g2_o21ai_1 _15147_ (.B1(_08479_),
    .Y(_01662_),
    .A1(net322),
    .A2(net473));
 sg13g2_nand2_1 _15148_ (.Y(_08480_),
    .A(\dp.rf.rf[25][3] ),
    .B(net473));
 sg13g2_o21ai_1 _15149_ (.B1(_08480_),
    .Y(_01663_),
    .A1(net318),
    .A2(net473));
 sg13g2_mux2_1 _15150_ (.A0(\dp.rf.rf[25][4] ),
    .A1(net290),
    .S(net477),
    .X(_01664_));
 sg13g2_nand2_1 _15151_ (.Y(_08481_),
    .A(\dp.rf.rf[25][5] ),
    .B(net471));
 sg13g2_o21ai_1 _15152_ (.B1(_08481_),
    .Y(_01665_),
    .A1(net312),
    .A2(net471));
 sg13g2_nand2_1 _15153_ (.Y(_08482_),
    .A(\dp.rf.rf[25][6] ),
    .B(net472));
 sg13g2_o21ai_1 _15154_ (.B1(_08482_),
    .Y(_01666_),
    .A1(net287),
    .A2(net472));
 sg13g2_nand2_1 _15155_ (.Y(_08483_),
    .A(\dp.rf.rf[25][7] ),
    .B(net472));
 sg13g2_o21ai_1 _15156_ (.B1(_08483_),
    .Y(_01667_),
    .A1(net284),
    .A2(net472));
 sg13g2_nand2_1 _15157_ (.Y(_08484_),
    .A(\dp.rf.rf[25][8] ),
    .B(net474));
 sg13g2_o21ai_1 _15158_ (.B1(_08484_),
    .Y(_01668_),
    .A1(net278),
    .A2(net474));
 sg13g2_buf_1 output112 (.A(net112),
    .X(pc[20]));
 sg13g2_nand2_1 _15160_ (.Y(_08486_),
    .A(\dp.rf.rf[25][9] ),
    .B(net471));
 sg13g2_o21ai_1 _15161_ (.B1(_08486_),
    .Y(_01669_),
    .A1(net271),
    .A2(net471));
 sg13g2_nand2_1 _15162_ (.Y(_08487_),
    .A(\dp.rf.rf[25][10] ),
    .B(net473));
 sg13g2_o21ai_1 _15163_ (.B1(_08487_),
    .Y(_01670_),
    .A1(net268),
    .A2(net473));
 sg13g2_nand2_1 _15164_ (.Y(_08488_),
    .A(\dp.rf.rf[25][11] ),
    .B(net474));
 sg13g2_o21ai_1 _15165_ (.B1(_08488_),
    .Y(_01671_),
    .A1(net262),
    .A2(net473));
 sg13g2_buf_1 output111 (.A(net111),
    .X(pc[1]));
 sg13g2_nand2_1 _15167_ (.Y(_08490_),
    .A(\dp.rf.rf[25][12] ),
    .B(net472));
 sg13g2_o21ai_1 _15168_ (.B1(_08490_),
    .Y(_01672_),
    .A1(net256),
    .A2(net472));
 sg13g2_mux2_1 _15169_ (.A0(\dp.rf.rf[25][13] ),
    .A1(net251),
    .S(net477),
    .X(_01673_));
 sg13g2_nor2_1 _15170_ (.A(\dp.rf.rf[25][14] ),
    .B(net477),
    .Y(_08491_));
 sg13g2_a21oi_1 _15171_ (.A1(net247),
    .A2(net477),
    .Y(_01674_),
    .B1(_08491_));
 sg13g2_nand2_1 _15172_ (.Y(_08492_),
    .A(\dp.rf.rf[25][15] ),
    .B(net471));
 sg13g2_o21ai_1 _15173_ (.B1(_08492_),
    .Y(_01675_),
    .A1(net240),
    .A2(net471));
 sg13g2_nand2_1 _15174_ (.Y(_08493_),
    .A(\dp.rf.rf[25][16] ),
    .B(net471));
 sg13g2_o21ai_1 _15175_ (.B1(_08493_),
    .Y(_01676_),
    .A1(net234),
    .A2(net471));
 sg13g2_nor2_1 _15176_ (.A(\dp.rf.rf[25][17] ),
    .B(net477),
    .Y(_08494_));
 sg13g2_a21oi_1 _15177_ (.A1(net231),
    .A2(net477),
    .Y(_01677_),
    .B1(_08494_));
 sg13g2_nand2_1 _15178_ (.Y(_08495_),
    .A(\dp.rf.rf[25][18] ),
    .B(net470));
 sg13g2_o21ai_1 _15179_ (.B1(_08495_),
    .Y(_01678_),
    .A1(net225),
    .A2(net470));
 sg13g2_nand2_1 _15180_ (.Y(_08496_),
    .A(\dp.rf.rf[25][19] ),
    .B(net470));
 sg13g2_o21ai_1 _15181_ (.B1(_08496_),
    .Y(_01679_),
    .A1(net220),
    .A2(net470));
 sg13g2_nor2_1 _15182_ (.A(\dp.rf.rf[25][20] ),
    .B(net476),
    .Y(_08497_));
 sg13g2_a21oi_1 _15183_ (.A1(net217),
    .A2(net476),
    .Y(_01680_),
    .B1(_08497_));
 sg13g2_nand2_1 _15184_ (.Y(_08498_),
    .A(\dp.rf.rf[25][21] ),
    .B(net469));
 sg13g2_o21ai_1 _15185_ (.B1(_08498_),
    .Y(_01681_),
    .A1(net211),
    .A2(net469));
 sg13g2_nor2_1 _15186_ (.A(\dp.rf.rf[25][22] ),
    .B(net476),
    .Y(_08499_));
 sg13g2_a21oi_1 _15187_ (.A1(_07639_),
    .A2(net476),
    .Y(_01682_),
    .B1(_08499_));
 sg13g2_nand2_1 _15188_ (.Y(_08500_),
    .A(\dp.rf.rf[25][23] ),
    .B(net468));
 sg13g2_o21ai_1 _15189_ (.B1(_08500_),
    .Y(_01683_),
    .A1(net201),
    .A2(net468));
 sg13g2_nand2_1 _15190_ (.Y(_08501_),
    .A(\dp.rf.rf[25][24] ),
    .B(net475));
 sg13g2_o21ai_1 _15191_ (.B1(_08501_),
    .Y(_01684_),
    .A1(net197),
    .A2(net475));
 sg13g2_nand2_1 _15192_ (.Y(_08502_),
    .A(\dp.rf.rf[25][25] ),
    .B(net468));
 sg13g2_o21ai_1 _15193_ (.B1(_08502_),
    .Y(_01685_),
    .A1(net193),
    .A2(net468));
 sg13g2_nand2_1 _15194_ (.Y(_08503_),
    .A(\dp.rf.rf[25][26] ),
    .B(net468));
 sg13g2_o21ai_1 _15195_ (.B1(_08503_),
    .Y(_01686_),
    .A1(net183),
    .A2(net468));
 sg13g2_nand2_1 _15196_ (.Y(_08504_),
    .A(\dp.rf.rf[25][27] ),
    .B(net468));
 sg13g2_o21ai_1 _15197_ (.B1(_08504_),
    .Y(_01687_),
    .A1(net179),
    .A2(net468));
 sg13g2_nand2_1 _15198_ (.Y(_08505_),
    .A(\dp.rf.rf[25][28] ),
    .B(net469));
 sg13g2_o21ai_1 _15199_ (.B1(_08505_),
    .Y(_01688_),
    .A1(net308),
    .A2(net469));
 sg13g2_nor2_1 _15200_ (.A(\dp.rf.rf[25][29] ),
    .B(net476),
    .Y(_08506_));
 sg13g2_a21oi_1 _15201_ (.A1(net175),
    .A2(net476),
    .Y(_01689_),
    .B1(_08506_));
 sg13g2_nor2_1 _15202_ (.A(\dp.rf.rf[25][30] ),
    .B(net476),
    .Y(_08507_));
 sg13g2_a21oi_1 _15203_ (.A1(net172),
    .A2(net476),
    .Y(_01690_),
    .B1(_08507_));
 sg13g2_nand2_1 _15204_ (.Y(_08508_),
    .A(\dp.rf.rf[25][31] ),
    .B(net470));
 sg13g2_o21ai_1 _15205_ (.B1(_08508_),
    .Y(_01691_),
    .A1(net165),
    .A2(net470));
 sg13g2_nor2_2 _15206_ (.A(_07924_),
    .B(_08468_),
    .Y(_08509_));
 sg13g2_buf_1 output110 (.A(net110),
    .X(pc[19]));
 sg13g2_nor2_1 _15208_ (.A(\dp.rf.rf[26][0] ),
    .B(_08509_),
    .Y(_08511_));
 sg13g2_a21oi_1 _15209_ (.A1(net303),
    .A2(_08509_),
    .Y(_01692_),
    .B1(_08511_));
 sg13g2_nand3_1 _15210_ (.B(_07745_),
    .C(_07930_),
    .A(net3),
    .Y(_08512_));
 sg13g2_buf_1 output109 (.A(net109),
    .X(pc[18]));
 sg13g2_buf_1 output108 (.A(net108),
    .X(pc[17]));
 sg13g2_buf_1 output107 (.A(net107),
    .X(pc[16]));
 sg13g2_nand2_1 _15214_ (.Y(_08516_),
    .A(\dp.rf.rf[26][1] ),
    .B(net706));
 sg13g2_o21ai_1 _15215_ (.B1(_08516_),
    .Y(_01693_),
    .A1(net298),
    .A2(net706));
 sg13g2_nand2_1 _15216_ (.Y(_02078_),
    .A(\dp.rf.rf[26][2] ),
    .B(net707));
 sg13g2_o21ai_1 _15217_ (.B1(_02078_),
    .Y(_01694_),
    .A1(net323),
    .A2(net707));
 sg13g2_nand2_1 _15218_ (.Y(_02079_),
    .A(\dp.rf.rf[26][3] ),
    .B(net706));
 sg13g2_o21ai_1 _15219_ (.B1(_02079_),
    .Y(_01695_),
    .A1(net318),
    .A2(net706));
 sg13g2_mux2_1 _15220_ (.A0(\dp.rf.rf[26][4] ),
    .A1(net290),
    .S(_08509_),
    .X(_01696_));
 sg13g2_buf_1 output106 (.A(net106),
    .X(pc[15]));
 sg13g2_nand2_1 _15222_ (.Y(_02081_),
    .A(\dp.rf.rf[26][5] ),
    .B(net705));
 sg13g2_o21ai_1 _15223_ (.B1(_02081_),
    .Y(_01697_),
    .A1(net312),
    .A2(net704));
 sg13g2_nand2_1 _15224_ (.Y(_02082_),
    .A(\dp.rf.rf[26][6] ),
    .B(net705));
 sg13g2_o21ai_1 _15225_ (.B1(_02082_),
    .Y(_01698_),
    .A1(net289),
    .A2(net705));
 sg13g2_nand2_1 _15226_ (.Y(_02083_),
    .A(\dp.rf.rf[26][7] ),
    .B(net705));
 sg13g2_o21ai_1 _15227_ (.B1(_02083_),
    .Y(_01699_),
    .A1(net283),
    .A2(net705));
 sg13g2_nand2_1 _15228_ (.Y(_02084_),
    .A(\dp.rf.rf[26][8] ),
    .B(net707));
 sg13g2_o21ai_1 _15229_ (.B1(_02084_),
    .Y(_01700_),
    .A1(net278),
    .A2(net707));
 sg13g2_nand2_1 _15230_ (.Y(_02085_),
    .A(\dp.rf.rf[26][9] ),
    .B(net704));
 sg13g2_o21ai_1 _15231_ (.B1(_02085_),
    .Y(_01701_),
    .A1(net271),
    .A2(net704));
 sg13g2_nand2_1 _15232_ (.Y(_02086_),
    .A(\dp.rf.rf[26][10] ),
    .B(net706));
 sg13g2_o21ai_1 _15233_ (.B1(_02086_),
    .Y(_01702_),
    .A1(net268),
    .A2(net706));
 sg13g2_nand2_1 _15234_ (.Y(_02087_),
    .A(\dp.rf.rf[26][11] ),
    .B(net706));
 sg13g2_o21ai_1 _15235_ (.B1(_02087_),
    .Y(_01703_),
    .A1(net262),
    .A2(net706));
 sg13g2_buf_1 output105 (.A(net105),
    .X(pc[14]));
 sg13g2_nand2_1 _15237_ (.Y(_02089_),
    .A(\dp.rf.rf[26][12] ),
    .B(net704));
 sg13g2_o21ai_1 _15238_ (.B1(_02089_),
    .Y(_01704_),
    .A1(net258),
    .A2(net705));
 sg13g2_mux2_1 _15239_ (.A0(\dp.rf.rf[26][13] ),
    .A1(net251),
    .S(_08509_),
    .X(_01705_));
 sg13g2_buf_1 output104 (.A(net104),
    .X(pc[13]));
 sg13g2_nand2_1 _15241_ (.Y(_02091_),
    .A(\dp.rf.rf[26][14] ),
    .B(net702));
 sg13g2_o21ai_1 _15242_ (.B1(_02091_),
    .Y(_01706_),
    .A1(net246),
    .A2(net702));
 sg13g2_nand2_1 _15243_ (.Y(_02092_),
    .A(\dp.rf.rf[26][15] ),
    .B(net704));
 sg13g2_o21ai_1 _15244_ (.B1(_02092_),
    .Y(_01707_),
    .A1(net242),
    .A2(net704));
 sg13g2_buf_1 output103 (.A(net103),
    .X(pc[12]));
 sg13g2_nand2_1 _15246_ (.Y(_02094_),
    .A(\dp.rf.rf[26][16] ),
    .B(net704));
 sg13g2_o21ai_1 _15247_ (.B1(_02094_),
    .Y(_01708_),
    .A1(net235),
    .A2(net704));
 sg13g2_nand2_1 _15248_ (.Y(_02095_),
    .A(\dp.rf.rf[26][17] ),
    .B(net708));
 sg13g2_o21ai_1 _15249_ (.B1(_02095_),
    .Y(_01709_),
    .A1(net231),
    .A2(net703));
 sg13g2_nand2_1 _15250_ (.Y(_02096_),
    .A(\dp.rf.rf[26][18] ),
    .B(net703));
 sg13g2_o21ai_1 _15251_ (.B1(_02096_),
    .Y(_01710_),
    .A1(net225),
    .A2(net703));
 sg13g2_nand2_1 _15252_ (.Y(_02097_),
    .A(\dp.rf.rf[26][19] ),
    .B(net702));
 sg13g2_o21ai_1 _15253_ (.B1(_02097_),
    .Y(_01711_),
    .A1(net219),
    .A2(net702));
 sg13g2_buf_1 output102 (.A(net102),
    .X(pc[11]));
 sg13g2_nand2_1 _15255_ (.Y(_02099_),
    .A(\dp.rf.rf[26][20] ),
    .B(net703));
 sg13g2_o21ai_1 _15256_ (.B1(_02099_),
    .Y(_01712_),
    .A1(net217),
    .A2(net703));
 sg13g2_nand2_1 _15257_ (.Y(_02100_),
    .A(\dp.rf.rf[26][21] ),
    .B(net701));
 sg13g2_o21ai_1 _15258_ (.B1(_02100_),
    .Y(_01713_),
    .A1(net211),
    .A2(net701));
 sg13g2_nor2_1 _15259_ (.A(\dp.rf.rf[26][22] ),
    .B(_08509_),
    .Y(_02101_));
 sg13g2_a21oi_1 _15260_ (.A1(net207),
    .A2(_08509_),
    .Y(_01714_),
    .B1(_02101_));
 sg13g2_nand2_1 _15261_ (.Y(_02102_),
    .A(\dp.rf.rf[26][23] ),
    .B(net700));
 sg13g2_o21ai_1 _15262_ (.B1(_02102_),
    .Y(_01715_),
    .A1(net200),
    .A2(net700));
 sg13g2_nand2_1 _15263_ (.Y(_02103_),
    .A(\dp.rf.rf[26][24] ),
    .B(net701));
 sg13g2_o21ai_1 _15264_ (.B1(_02103_),
    .Y(_01716_),
    .A1(net197),
    .A2(net701));
 sg13g2_nand2_1 _15265_ (.Y(_02104_),
    .A(\dp.rf.rf[26][25] ),
    .B(net700));
 sg13g2_o21ai_1 _15266_ (.B1(_02104_),
    .Y(_01717_),
    .A1(net190),
    .A2(net700));
 sg13g2_nand2_1 _15267_ (.Y(_02105_),
    .A(\dp.rf.rf[26][26] ),
    .B(net700));
 sg13g2_o21ai_1 _15268_ (.B1(_02105_),
    .Y(_01718_),
    .A1(net183),
    .A2(net700));
 sg13g2_nand2_1 _15269_ (.Y(_02106_),
    .A(\dp.rf.rf[26][27] ),
    .B(net700));
 sg13g2_o21ai_1 _15270_ (.B1(_02106_),
    .Y(_01719_),
    .A1(net179),
    .A2(net700));
 sg13g2_nand2_1 _15271_ (.Y(_02107_),
    .A(\dp.rf.rf[26][28] ),
    .B(net701));
 sg13g2_o21ai_1 _15272_ (.B1(_02107_),
    .Y(_01720_),
    .A1(net308),
    .A2(net701));
 sg13g2_nor2_1 _15273_ (.A(\dp.rf.rf[26][29] ),
    .B(_08509_),
    .Y(_02108_));
 sg13g2_a21oi_1 _15274_ (.A1(net175),
    .A2(_08509_),
    .Y(_01721_),
    .B1(_02108_));
 sg13g2_nand2_1 _15275_ (.Y(_02109_),
    .A(\dp.rf.rf[26][30] ),
    .B(net703));
 sg13g2_o21ai_1 _15276_ (.B1(_02109_),
    .Y(_01722_),
    .A1(net172),
    .A2(net703));
 sg13g2_nand2_1 _15277_ (.Y(_02110_),
    .A(\dp.rf.rf[26][31] ),
    .B(net702));
 sg13g2_o21ai_1 _15278_ (.B1(_02110_),
    .Y(_01723_),
    .A1(net166),
    .A2(net702));
 sg13g2_nand2b_1 _15279_ (.Y(_02111_),
    .B(_07841_),
    .A_N(_07787_));
 sg13g2_buf_1 output101 (.A(net101),
    .X(pc[10]));
 sg13g2_buf_1 output100 (.A(net100),
    .X(pc[0]));
 sg13g2_buf_1 output99 (.A(net99),
    .X(memwrite));
 sg13g2_nand2_1 _15283_ (.Y(_02115_),
    .A(\dp.rf.rf[28][0] ),
    .B(net693));
 sg13g2_o21ai_1 _15284_ (.B1(_02115_),
    .Y(_01724_),
    .A1(net302),
    .A2(net693));
 sg13g2_buf_1 output98 (.A(net829),
    .X(memread));
 sg13g2_nand2_1 _15286_ (.Y(_02117_),
    .A(\dp.rf.rf[28][1] ),
    .B(net697));
 sg13g2_o21ai_1 _15287_ (.B1(_02117_),
    .Y(_01725_),
    .A1(net299),
    .A2(net697));
 sg13g2_buf_1 output97 (.A(net97),
    .X(aluout[9]));
 sg13g2_nand2_1 _15289_ (.Y(_02119_),
    .A(\dp.rf.rf[28][2] ),
    .B(net697));
 sg13g2_o21ai_1 _15290_ (.B1(_02119_),
    .Y(_01726_),
    .A1(net322),
    .A2(net697));
 sg13g2_buf_1 output96 (.A(net96),
    .X(aluout[8]));
 sg13g2_nand2_1 _15292_ (.Y(_02121_),
    .A(\dp.rf.rf[28][3] ),
    .B(net698));
 sg13g2_o21ai_1 _15293_ (.B1(_02121_),
    .Y(_01727_),
    .A1(net318),
    .A2(net698));
 sg13g2_nor2_2 _15294_ (.A(_07787_),
    .B(_08016_),
    .Y(_02122_));
 sg13g2_buf_1 output95 (.A(net95),
    .X(aluout[7]));
 sg13g2_mux2_1 _15296_ (.A0(\dp.rf.rf[28][4] ),
    .A1(net292),
    .S(_02122_),
    .X(_01728_));
 sg13g2_buf_1 output94 (.A(net94),
    .X(aluout[6]));
 sg13g2_buf_1 output93 (.A(net93),
    .X(aluout[5]));
 sg13g2_nand2_1 _15299_ (.Y(_02126_),
    .A(\dp.rf.rf[28][5] ),
    .B(net695));
 sg13g2_o21ai_1 _15300_ (.B1(_02126_),
    .Y(_01729_),
    .A1(net312),
    .A2(net695));
 sg13g2_buf_1 output92 (.A(net92),
    .X(aluout[4]));
 sg13g2_nand2_1 _15302_ (.Y(_02128_),
    .A(\dp.rf.rf[28][6] ),
    .B(net695));
 sg13g2_o21ai_1 _15303_ (.B1(_02128_),
    .Y(_01730_),
    .A1(net287),
    .A2(net695));
 sg13g2_buf_1 output91 (.A(net91),
    .X(aluout[3]));
 sg13g2_nand2_1 _15305_ (.Y(_02130_),
    .A(\dp.rf.rf[28][7] ),
    .B(net696));
 sg13g2_o21ai_1 _15306_ (.B1(_02130_),
    .Y(_01731_),
    .A1(net284),
    .A2(net696));
 sg13g2_buf_1 output90 (.A(net90),
    .X(aluout[31]));
 sg13g2_nand2_1 _15308_ (.Y(_02132_),
    .A(\dp.rf.rf[28][8] ),
    .B(net698));
 sg13g2_o21ai_1 _15309_ (.B1(_02132_),
    .Y(_01732_),
    .A1(net279),
    .A2(net698));
 sg13g2_buf_1 output89 (.A(net89),
    .X(aluout[30]));
 sg13g2_nand2_1 _15311_ (.Y(_02134_),
    .A(\dp.rf.rf[28][9] ),
    .B(net696));
 sg13g2_o21ai_1 _15312_ (.B1(_02134_),
    .Y(_01733_),
    .A1(net272),
    .A2(net696));
 sg13g2_buf_1 output88 (.A(net88),
    .X(aluout[2]));
 sg13g2_nand2_1 _15314_ (.Y(_02136_),
    .A(\dp.rf.rf[28][10] ),
    .B(net697));
 sg13g2_o21ai_1 _15315_ (.B1(_02136_),
    .Y(_01734_),
    .A1(net268),
    .A2(net697));
 sg13g2_buf_1 output87 (.A(net87),
    .X(aluout[29]));
 sg13g2_buf_1 output86 (.A(net86),
    .X(aluout[28]));
 sg13g2_nand2_1 _15318_ (.Y(_02139_),
    .A(\dp.rf.rf[28][11] ),
    .B(net697));
 sg13g2_o21ai_1 _15319_ (.B1(_02139_),
    .Y(_01735_),
    .A1(net262),
    .A2(net697));
 sg13g2_buf_1 output85 (.A(net85),
    .X(aluout[27]));
 sg13g2_nand2_1 _15321_ (.Y(_02141_),
    .A(\dp.rf.rf[28][12] ),
    .B(net695));
 sg13g2_o21ai_1 _15322_ (.B1(_02141_),
    .Y(_01736_),
    .A1(net256),
    .A2(net695));
 sg13g2_mux2_1 _15323_ (.A0(\dp.rf.rf[28][13] ),
    .A1(net251),
    .S(_02122_),
    .X(_01737_));
 sg13g2_nand2_1 _15324_ (.Y(_02142_),
    .A(\dp.rf.rf[28][14] ),
    .B(net694));
 sg13g2_o21ai_1 _15325_ (.B1(_02142_),
    .Y(_01738_),
    .A1(net248),
    .A2(net699));
 sg13g2_buf_1 output84 (.A(net84),
    .X(aluout[26]));
 sg13g2_nand2_1 _15327_ (.Y(_02144_),
    .A(\dp.rf.rf[28][15] ),
    .B(net695));
 sg13g2_o21ai_1 _15328_ (.B1(_02144_),
    .Y(_01739_),
    .A1(net241),
    .A2(net695));
 sg13g2_buf_1 output83 (.A(net83),
    .X(aluout[25]));
 sg13g2_buf_1 output82 (.A(net82),
    .X(aluout[24]));
 sg13g2_nand2_1 _15331_ (.Y(_02147_),
    .A(\dp.rf.rf[28][16] ),
    .B(net696));
 sg13g2_o21ai_1 _15332_ (.B1(_02147_),
    .Y(_01740_),
    .A1(net234),
    .A2(net696));
 sg13g2_nor2_1 _15333_ (.A(\dp.rf.rf[28][17] ),
    .B(net690),
    .Y(_02148_));
 sg13g2_a21oi_1 _15334_ (.A1(net231),
    .A2(net690),
    .Y(_01741_),
    .B1(_02148_));
 sg13g2_buf_1 output81 (.A(net81),
    .X(aluout[23]));
 sg13g2_nand2_1 _15336_ (.Y(_02150_),
    .A(\dp.rf.rf[28][18] ),
    .B(net694));
 sg13g2_o21ai_1 _15337_ (.B1(_02150_),
    .Y(_01742_),
    .A1(net226),
    .A2(net694));
 sg13g2_buf_1 output80 (.A(net80),
    .X(aluout[22]));
 sg13g2_nand2_1 _15339_ (.Y(_02152_),
    .A(\dp.rf.rf[28][19] ),
    .B(net693));
 sg13g2_o21ai_1 _15340_ (.B1(_02152_),
    .Y(_01743_),
    .A1(net221),
    .A2(net693));
 sg13g2_nand2_1 _15341_ (.Y(_02153_),
    .A(\dp.rf.rf[28][20] ),
    .B(net694));
 sg13g2_o21ai_1 _15342_ (.B1(_02153_),
    .Y(_01744_),
    .A1(net216),
    .A2(net694));
 sg13g2_buf_1 output79 (.A(net79),
    .X(aluout[21]));
 sg13g2_nand2_1 _15344_ (.Y(_02155_),
    .A(\dp.rf.rf[28][21] ),
    .B(net692));
 sg13g2_o21ai_1 _15345_ (.B1(_02155_),
    .Y(_01745_),
    .A1(net212),
    .A2(net692));
 sg13g2_nor2_1 _15346_ (.A(\dp.rf.rf[28][22] ),
    .B(net690),
    .Y(_02156_));
 sg13g2_a21oi_1 _15347_ (.A1(net207),
    .A2(net690),
    .Y(_01746_),
    .B1(_02156_));
 sg13g2_buf_1 output78 (.A(net78),
    .X(aluout[20]));
 sg13g2_nand2_1 _15349_ (.Y(_02158_),
    .A(\dp.rf.rf[28][23] ),
    .B(net691));
 sg13g2_o21ai_1 _15350_ (.B1(_02158_),
    .Y(_01747_),
    .A1(net200),
    .A2(net691));
 sg13g2_buf_1 output77 (.A(net77),
    .X(aluout[1]));
 sg13g2_nand2_1 _15352_ (.Y(_02160_),
    .A(\dp.rf.rf[28][24] ),
    .B(net694));
 sg13g2_o21ai_1 _15353_ (.B1(_02160_),
    .Y(_01748_),
    .A1(net198),
    .A2(net694));
 sg13g2_buf_1 output76 (.A(net76),
    .X(aluout[19]));
 sg13g2_nand2_1 _15355_ (.Y(_02162_),
    .A(\dp.rf.rf[28][25] ),
    .B(net691));
 sg13g2_o21ai_1 _15356_ (.B1(_02162_),
    .Y(_01749_),
    .A1(net189),
    .A2(net691));
 sg13g2_buf_1 output75 (.A(net75),
    .X(aluout[18]));
 sg13g2_nand2_1 _15358_ (.Y(_02164_),
    .A(\dp.rf.rf[28][26] ),
    .B(net691));
 sg13g2_o21ai_1 _15359_ (.B1(_02164_),
    .Y(_01750_),
    .A1(net184),
    .A2(net691));
 sg13g2_buf_1 output74 (.A(net74),
    .X(aluout[17]));
 sg13g2_nand2_1 _15361_ (.Y(_02166_),
    .A(\dp.rf.rf[28][27] ),
    .B(net691));
 sg13g2_o21ai_1 _15362_ (.B1(_02166_),
    .Y(_01751_),
    .A1(net179),
    .A2(net691));
 sg13g2_buf_1 output73 (.A(net73),
    .X(aluout[16]));
 sg13g2_nand2_1 _15364_ (.Y(_02168_),
    .A(\dp.rf.rf[28][28] ),
    .B(net692));
 sg13g2_o21ai_1 _15365_ (.B1(_02168_),
    .Y(_01752_),
    .A1(net306),
    .A2(net692));
 sg13g2_nor2_1 _15366_ (.A(\dp.rf.rf[28][29] ),
    .B(net690),
    .Y(_02169_));
 sg13g2_a21oi_1 _15367_ (.A1(net174),
    .A2(net690),
    .Y(_01753_),
    .B1(_02169_));
 sg13g2_nor2_1 _15368_ (.A(\dp.rf.rf[28][30] ),
    .B(net690),
    .Y(_02170_));
 sg13g2_a21oi_1 _15369_ (.A1(net173),
    .A2(net690),
    .Y(_01754_),
    .B1(_02170_));
 sg13g2_buf_1 output72 (.A(net72),
    .X(aluout[15]));
 sg13g2_nand2_1 _15371_ (.Y(_02172_),
    .A(\dp.rf.rf[28][31] ),
    .B(net693));
 sg13g2_o21ai_1 _15372_ (.B1(_02172_),
    .Y(_01755_),
    .A1(net166),
    .A2(net693));
 sg13g2_nand2_1 _15373_ (.Y(_02173_),
    .A(net1245),
    .B(_07395_));
 sg13g2_or2_1 _15374_ (.X(_02174_),
    .B(_08468_),
    .A(_02173_));
 sg13g2_buf_1 output71 (.A(net71),
    .X(aluout[14]));
 sg13g2_buf_1 output70 (.A(net70),
    .X(aluout[13]));
 sg13g2_buf_1 output69 (.A(net69),
    .X(aluout[12]));
 sg13g2_nand2_1 _15378_ (.Y(_02178_),
    .A(\dp.rf.rf[27][0] ),
    .B(net463));
 sg13g2_o21ai_1 _15379_ (.B1(_02178_),
    .Y(_01756_),
    .A1(net303),
    .A2(net463));
 sg13g2_nand2_1 _15380_ (.Y(_02179_),
    .A(\dp.rf.rf[27][1] ),
    .B(net465));
 sg13g2_o21ai_1 _15381_ (.B1(_02179_),
    .Y(_01757_),
    .A1(net298),
    .A2(net465));
 sg13g2_nand2_1 _15382_ (.Y(_02180_),
    .A(\dp.rf.rf[27][2] ),
    .B(net466));
 sg13g2_o21ai_1 _15383_ (.B1(_02180_),
    .Y(_01758_),
    .A1(net323),
    .A2(net466));
 sg13g2_nand2_1 _15384_ (.Y(_02181_),
    .A(\dp.rf.rf[27][3] ),
    .B(net465));
 sg13g2_o21ai_1 _15385_ (.B1(_02181_),
    .Y(_01759_),
    .A1(net318),
    .A2(net465));
 sg13g2_mux2_1 _15386_ (.A0(net292),
    .A1(\dp.rf.rf[27][4] ),
    .S(net461),
    .X(_01760_));
 sg13g2_nand2_1 _15387_ (.Y(_02182_),
    .A(\dp.rf.rf[27][5] ),
    .B(net464));
 sg13g2_o21ai_1 _15388_ (.B1(_02182_),
    .Y(_01761_),
    .A1(net312),
    .A2(net464));
 sg13g2_nand2_1 _15389_ (.Y(_02183_),
    .A(\dp.rf.rf[27][6] ),
    .B(net464));
 sg13g2_o21ai_1 _15390_ (.B1(_02183_),
    .Y(_01762_),
    .A1(net288),
    .A2(net464));
 sg13g2_nand2_1 _15391_ (.Y(_02184_),
    .A(\dp.rf.rf[27][7] ),
    .B(net464));
 sg13g2_o21ai_1 _15392_ (.B1(_02184_),
    .Y(_01763_),
    .A1(net283),
    .A2(net464));
 sg13g2_nand2_1 _15393_ (.Y(_02185_),
    .A(\dp.rf.rf[27][8] ),
    .B(net466));
 sg13g2_o21ai_1 _15394_ (.B1(_02185_),
    .Y(_01764_),
    .A1(net278),
    .A2(net466));
 sg13g2_buf_1 output68 (.A(net68),
    .X(aluout[11]));
 sg13g2_nand2_1 _15396_ (.Y(_02187_),
    .A(\dp.rf.rf[27][9] ),
    .B(net463));
 sg13g2_o21ai_1 _15397_ (.B1(_02187_),
    .Y(_01765_),
    .A1(net271),
    .A2(net463));
 sg13g2_nand2_1 _15398_ (.Y(_02188_),
    .A(\dp.rf.rf[27][10] ),
    .B(net465));
 sg13g2_o21ai_1 _15399_ (.B1(_02188_),
    .Y(_01766_),
    .A1(net269),
    .A2(net465));
 sg13g2_buf_1 output67 (.A(net67),
    .X(aluout[10]));
 sg13g2_nand2_1 _15401_ (.Y(_02190_),
    .A(\dp.rf.rf[27][11] ),
    .B(net465));
 sg13g2_o21ai_1 _15402_ (.B1(_02190_),
    .Y(_01767_),
    .A1(net262),
    .A2(net465));
 sg13g2_nand2_1 _15403_ (.Y(_02191_),
    .A(\dp.rf.rf[27][12] ),
    .B(net464));
 sg13g2_o21ai_1 _15404_ (.B1(_02191_),
    .Y(_01768_),
    .A1(net256),
    .A2(net464));
 sg13g2_mux2_1 _15405_ (.A0(net251),
    .A1(\dp.rf.rf[27][13] ),
    .S(net461),
    .X(_01769_));
 sg13g2_nand2_1 _15406_ (.Y(_02192_),
    .A(\dp.rf.rf[27][14] ),
    .B(net459));
 sg13g2_o21ai_1 _15407_ (.B1(_02192_),
    .Y(_01770_),
    .A1(net247),
    .A2(net459));
 sg13g2_nand2_1 _15408_ (.Y(_02193_),
    .A(\dp.rf.rf[27][15] ),
    .B(net463));
 sg13g2_o21ai_1 _15409_ (.B1(_02193_),
    .Y(_01771_),
    .A1(net242),
    .A2(net463));
 sg13g2_nand2_1 _15410_ (.Y(_02194_),
    .A(\dp.rf.rf[27][16] ),
    .B(net463));
 sg13g2_o21ai_1 _15411_ (.B1(_02194_),
    .Y(_01772_),
    .A1(net235),
    .A2(net463));
 sg13g2_nand2_1 _15412_ (.Y(_02195_),
    .A(\dp.rf.rf[27][17] ),
    .B(net460));
 sg13g2_o21ai_1 _15413_ (.B1(_02195_),
    .Y(_01773_),
    .A1(net231),
    .A2(net460));
 sg13g2_nand2_1 _15414_ (.Y(_02196_),
    .A(\dp.rf.rf[27][18] ),
    .B(net462));
 sg13g2_o21ai_1 _15415_ (.B1(_02196_),
    .Y(_01774_),
    .A1(net224),
    .A2(net462));
 sg13g2_nand2_1 _15416_ (.Y(_02197_),
    .A(\dp.rf.rf[27][19] ),
    .B(net459));
 sg13g2_o21ai_1 _15417_ (.B1(_02197_),
    .Y(_01775_),
    .A1(net220),
    .A2(net459));
 sg13g2_buf_1 output66 (.A(net66),
    .X(aluout[0]));
 sg13g2_nand2_1 _15419_ (.Y(_02199_),
    .A(\dp.rf.rf[27][20] ),
    .B(net460));
 sg13g2_o21ai_1 _15420_ (.B1(_02199_),
    .Y(_01776_),
    .A1(net217),
    .A2(net460));
 sg13g2_nand2_1 _15421_ (.Y(_02200_),
    .A(\dp.rf.rf[27][21] ),
    .B(net458));
 sg13g2_o21ai_1 _15422_ (.B1(_02200_),
    .Y(_01777_),
    .A1(net211),
    .A2(net458));
 sg13g2_buf_1 input65 (.A(reset),
    .X(net65));
 sg13g2_nand2_1 _15424_ (.Y(_02202_),
    .A(\dp.rf.rf[27][22] ),
    .B(net460));
 sg13g2_o21ai_1 _15425_ (.B1(_02202_),
    .Y(_01778_),
    .A1(net207),
    .A2(net461));
 sg13g2_nand2_1 _15426_ (.Y(_02203_),
    .A(\dp.rf.rf[27][23] ),
    .B(net457));
 sg13g2_o21ai_1 _15427_ (.B1(_02203_),
    .Y(_01779_),
    .A1(net201),
    .A2(net457));
 sg13g2_nand2_1 _15428_ (.Y(_02204_),
    .A(\dp.rf.rf[27][24] ),
    .B(net458));
 sg13g2_o21ai_1 _15429_ (.B1(_02204_),
    .Y(_01780_),
    .A1(net197),
    .A2(net458));
 sg13g2_nand2_1 _15430_ (.Y(_02205_),
    .A(\dp.rf.rf[27][25] ),
    .B(net457));
 sg13g2_o21ai_1 _15431_ (.B1(_02205_),
    .Y(_01781_),
    .A1(net193),
    .A2(net457));
 sg13g2_nand2_1 _15432_ (.Y(_02206_),
    .A(\dp.rf.rf[27][26] ),
    .B(net457));
 sg13g2_o21ai_1 _15433_ (.B1(_02206_),
    .Y(_01782_),
    .A1(net183),
    .A2(net457));
 sg13g2_nand2_1 _15434_ (.Y(_02207_),
    .A(\dp.rf.rf[27][27] ),
    .B(net457));
 sg13g2_o21ai_1 _15435_ (.B1(_02207_),
    .Y(_01783_),
    .A1(net180),
    .A2(net457));
 sg13g2_nand2_1 _15436_ (.Y(_02208_),
    .A(\dp.rf.rf[27][28] ),
    .B(net458));
 sg13g2_o21ai_1 _15437_ (.B1(_02208_),
    .Y(_01784_),
    .A1(net308),
    .A2(net458));
 sg13g2_nand2_1 _15438_ (.Y(_02209_),
    .A(\dp.rf.rf[27][29] ),
    .B(net460));
 sg13g2_o21ai_1 _15439_ (.B1(_02209_),
    .Y(_01785_),
    .A1(net175),
    .A2(net460));
 sg13g2_nand2_1 _15440_ (.Y(_02210_),
    .A(\dp.rf.rf[27][30] ),
    .B(net460));
 sg13g2_o21ai_1 _15441_ (.B1(_02210_),
    .Y(_01786_),
    .A1(net172),
    .A2(net461));
 sg13g2_nand2_1 _15442_ (.Y(_02211_),
    .A(\dp.rf.rf[27][31] ),
    .B(net459));
 sg13g2_o21ai_1 _15443_ (.B1(_02211_),
    .Y(_01787_),
    .A1(net166),
    .A2(net459));
 sg13g2_nand2_1 _15444_ (.Y(_02212_),
    .A(_07840_),
    .B(_07930_));
 sg13g2_buf_1 input64 (.A(readdata[9]),
    .X(net64));
 sg13g2_buf_1 input63 (.A(readdata[8]),
    .X(net63));
 sg13g2_buf_1 input62 (.A(readdata[7]),
    .X(net62));
 sg13g2_nand2_1 _15448_ (.Y(_02216_),
    .A(\dp.rf.rf[2][0] ),
    .B(net684));
 sg13g2_o21ai_1 _15449_ (.B1(_02216_),
    .Y(_01788_),
    .A1(net300),
    .A2(net684));
 sg13g2_nand2_1 _15450_ (.Y(_02217_),
    .A(\dp.rf.rf[2][1] ),
    .B(net688));
 sg13g2_o21ai_1 _15451_ (.B1(_02217_),
    .Y(_01789_),
    .A1(net296),
    .A2(net688));
 sg13g2_nand2_1 _15452_ (.Y(_02218_),
    .A(\dp.rf.rf[2][2] ),
    .B(net688));
 sg13g2_o21ai_1 _15453_ (.B1(_02218_),
    .Y(_01790_),
    .A1(net321),
    .A2(net688));
 sg13g2_nand2_1 _15454_ (.Y(_02219_),
    .A(\dp.rf.rf[2][3] ),
    .B(net688));
 sg13g2_o21ai_1 _15455_ (.B1(_02219_),
    .Y(_01791_),
    .A1(net315),
    .A2(net688));
 sg13g2_mux2_1 _15456_ (.A0(net294),
    .A1(\dp.rf.rf[2][4] ),
    .S(net687),
    .X(_01792_));
 sg13g2_nand2_1 _15457_ (.Y(_02220_),
    .A(\dp.rf.rf[2][5] ),
    .B(net686));
 sg13g2_o21ai_1 _15458_ (.B1(_02220_),
    .Y(_01793_),
    .A1(net311),
    .A2(net686));
 sg13g2_nand2_1 _15459_ (.Y(_02221_),
    .A(\dp.rf.rf[2][6] ),
    .B(net685));
 sg13g2_o21ai_1 _15460_ (.B1(_02221_),
    .Y(_01794_),
    .A1(net286),
    .A2(net685));
 sg13g2_nand2_1 _15461_ (.Y(_02222_),
    .A(\dp.rf.rf[2][7] ),
    .B(net686));
 sg13g2_o21ai_1 _15462_ (.B1(_02222_),
    .Y(_01795_),
    .A1(net281),
    .A2(net686));
 sg13g2_nand2_1 _15463_ (.Y(_02223_),
    .A(\dp.rf.rf[2][8] ),
    .B(net689));
 sg13g2_o21ai_1 _15464_ (.B1(_02223_),
    .Y(_01796_),
    .A1(net277),
    .A2(net689));
 sg13g2_buf_1 input61 (.A(readdata[6]),
    .X(net61));
 sg13g2_nand2_1 _15466_ (.Y(_02225_),
    .A(\dp.rf.rf[2][9] ),
    .B(net684));
 sg13g2_o21ai_1 _15467_ (.B1(_02225_),
    .Y(_01797_),
    .A1(net274),
    .A2(net684));
 sg13g2_nand2_1 _15468_ (.Y(_02226_),
    .A(\dp.rf.rf[2][10] ),
    .B(net685));
 sg13g2_o21ai_1 _15469_ (.B1(_02226_),
    .Y(_01798_),
    .A1(net267),
    .A2(net685));
 sg13g2_buf_1 input60 (.A(readdata[5]),
    .X(net60));
 sg13g2_nand2_1 _15471_ (.Y(_02228_),
    .A(\dp.rf.rf[2][11] ),
    .B(net689));
 sg13g2_o21ai_1 _15472_ (.B1(_02228_),
    .Y(_01799_),
    .A1(net260),
    .A2(net689));
 sg13g2_nand2_1 _15473_ (.Y(_02229_),
    .A(\dp.rf.rf[2][12] ),
    .B(net688));
 sg13g2_o21ai_1 _15474_ (.B1(_02229_),
    .Y(_01800_),
    .A1(net254),
    .A2(net688));
 sg13g2_mux2_1 _15475_ (.A0(net253),
    .A1(\dp.rf.rf[2][13] ),
    .S(net689),
    .X(_01801_));
 sg13g2_nand2_1 _15476_ (.Y(_02230_),
    .A(\dp.rf.rf[2][14] ),
    .B(net679));
 sg13g2_o21ai_1 _15477_ (.B1(_02230_),
    .Y(_01802_),
    .A1(net247),
    .A2(net679));
 sg13g2_nand2_1 _15478_ (.Y(_02231_),
    .A(\dp.rf.rf[2][15] ),
    .B(net685));
 sg13g2_o21ai_1 _15479_ (.B1(_02231_),
    .Y(_01803_),
    .A1(net244),
    .A2(net685));
 sg13g2_nand2_1 _15480_ (.Y(_02232_),
    .A(\dp.rf.rf[2][16] ),
    .B(net685));
 sg13g2_o21ai_1 _15481_ (.B1(_02232_),
    .Y(_01804_),
    .A1(net237),
    .A2(net685));
 sg13g2_nand2_1 _15482_ (.Y(_02233_),
    .A(\dp.rf.rf[2][17] ),
    .B(net680));
 sg13g2_o21ai_1 _15483_ (.B1(_02233_),
    .Y(_01805_),
    .A1(net229),
    .A2(net683));
 sg13g2_nand2_1 _15484_ (.Y(_02234_),
    .A(\dp.rf.rf[2][18] ),
    .B(net684));
 sg13g2_o21ai_1 _15485_ (.B1(_02234_),
    .Y(_01806_),
    .A1(net228),
    .A2(net684));
 sg13g2_nand2_1 _15486_ (.Y(_02235_),
    .A(\dp.rf.rf[2][19] ),
    .B(net684));
 sg13g2_o21ai_1 _15487_ (.B1(_02235_),
    .Y(_01807_),
    .A1(net222),
    .A2(net684));
 sg13g2_buf_1 input59 (.A(readdata[4]),
    .X(net59));
 sg13g2_nand2_1 _15489_ (.Y(_02237_),
    .A(\dp.rf.rf[2][20] ),
    .B(net681));
 sg13g2_o21ai_1 _15490_ (.B1(_02237_),
    .Y(_01808_),
    .A1(net215),
    .A2(net681));
 sg13g2_nand2_1 _15491_ (.Y(_02238_),
    .A(\dp.rf.rf[2][21] ),
    .B(net680));
 sg13g2_o21ai_1 _15492_ (.B1(_02238_),
    .Y(_01809_),
    .A1(net213),
    .A2(net680));
 sg13g2_buf_1 input58 (.A(readdata[3]),
    .X(net58));
 sg13g2_nand2_1 _15494_ (.Y(_02240_),
    .A(\dp.rf.rf[2][22] ),
    .B(net682));
 sg13g2_o21ai_1 _15495_ (.B1(_02240_),
    .Y(_01810_),
    .A1(net206),
    .A2(net682));
 sg13g2_nand2_1 _15496_ (.Y(_02241_),
    .A(\dp.rf.rf[2][23] ),
    .B(net679));
 sg13g2_o21ai_1 _15497_ (.B1(_02241_),
    .Y(_01811_),
    .A1(net203),
    .A2(net679));
 sg13g2_nand2_1 _15498_ (.Y(_02242_),
    .A(\dp.rf.rf[2][24] ),
    .B(net681));
 sg13g2_o21ai_1 _15499_ (.B1(_02242_),
    .Y(_01812_),
    .A1(net196),
    .A2(net681));
 sg13g2_nand2_1 _15500_ (.Y(_02243_),
    .A(\dp.rf.rf[2][25] ),
    .B(net680));
 sg13g2_o21ai_1 _15501_ (.B1(_02243_),
    .Y(_01813_),
    .A1(net192),
    .A2(net680));
 sg13g2_nand2_1 _15502_ (.Y(_02244_),
    .A(\dp.rf.rf[2][26] ),
    .B(net681));
 sg13g2_o21ai_1 _15503_ (.B1(_02244_),
    .Y(_01814_),
    .A1(net188),
    .A2(net681));
 sg13g2_nand2_1 _15504_ (.Y(_02245_),
    .A(\dp.rf.rf[2][27] ),
    .B(net679));
 sg13g2_o21ai_1 _15505_ (.B1(_02245_),
    .Y(_01815_),
    .A1(net181),
    .A2(net679));
 sg13g2_nand2_1 _15506_ (.Y(_02246_),
    .A(\dp.rf.rf[2][28] ),
    .B(net680));
 sg13g2_o21ai_1 _15507_ (.B1(_02246_),
    .Y(_01816_),
    .A1(net307),
    .A2(net680));
 sg13g2_nand2_1 _15508_ (.Y(_02247_),
    .A(\dp.rf.rf[2][29] ),
    .B(net681));
 sg13g2_o21ai_1 _15509_ (.B1(_02247_),
    .Y(_01817_),
    .A1(net177),
    .A2(net682));
 sg13g2_nand2_1 _15510_ (.Y(_02248_),
    .A(\dp.rf.rf[2][30] ),
    .B(net681));
 sg13g2_o21ai_1 _15511_ (.B1(_02248_),
    .Y(_01818_),
    .A1(net171),
    .A2(net682));
 sg13g2_nand2_1 _15512_ (.Y(_02249_),
    .A(\dp.rf.rf[2][31] ),
    .B(net679));
 sg13g2_o21ai_1 _15513_ (.B1(_02249_),
    .Y(_01819_),
    .A1(net168),
    .A2(net679));
 sg13g2_nand2b_2 _15514_ (.Y(_02250_),
    .B(_07930_),
    .A_N(_07787_));
 sg13g2_buf_1 input57 (.A(readdata[31]),
    .X(net57));
 sg13g2_buf_1 input56 (.A(readdata[30]),
    .X(net56));
 sg13g2_buf_1 input55 (.A(readdata[2]),
    .X(net55));
 sg13g2_buf_1 input54 (.A(readdata[29]),
    .X(net54));
 sg13g2_nand2_1 _15519_ (.Y(_02255_),
    .A(\dp.rf.rf[30][0] ),
    .B(net672));
 sg13g2_o21ai_1 _15520_ (.B1(_02255_),
    .Y(_01820_),
    .A1(net301),
    .A2(net672));
 sg13g2_nand2_1 _15521_ (.Y(_02256_),
    .A(\dp.rf.rf[30][1] ),
    .B(net677));
 sg13g2_o21ai_1 _15522_ (.B1(_02256_),
    .Y(_01821_),
    .A1(net298),
    .A2(net677));
 sg13g2_buf_1 input53 (.A(readdata[28]),
    .X(net53));
 sg13g2_nand2_1 _15524_ (.Y(_02258_),
    .A(\dp.rf.rf[30][2] ),
    .B(net678));
 sg13g2_o21ai_1 _15525_ (.B1(_02258_),
    .Y(_01822_),
    .A1(net322),
    .A2(net677));
 sg13g2_nand2_1 _15526_ (.Y(_02259_),
    .A(\dp.rf.rf[30][3] ),
    .B(net677));
 sg13g2_o21ai_1 _15527_ (.B1(_02259_),
    .Y(_01823_),
    .A1(net318),
    .A2(net677));
 sg13g2_nor2_2 _15528_ (.A(_07787_),
    .B(_07924_),
    .Y(_02260_));
 sg13g2_buf_1 input52 (.A(readdata[27]),
    .X(net52));
 sg13g2_mux2_1 _15530_ (.A0(\dp.rf.rf[30][4] ),
    .A1(net292),
    .S(_02260_),
    .X(_01824_));
 sg13g2_nand2_1 _15531_ (.Y(_02262_),
    .A(\dp.rf.rf[30][5] ),
    .B(net675));
 sg13g2_o21ai_1 _15532_ (.B1(_02262_),
    .Y(_01825_),
    .A1(net312),
    .A2(net675));
 sg13g2_nand2_1 _15533_ (.Y(_02263_),
    .A(\dp.rf.rf[30][6] ),
    .B(net675));
 sg13g2_o21ai_1 _15534_ (.B1(_02263_),
    .Y(_01826_),
    .A1(net287),
    .A2(net675));
 sg13g2_nand2_1 _15535_ (.Y(_02264_),
    .A(\dp.rf.rf[30][7] ),
    .B(net676));
 sg13g2_o21ai_1 _15536_ (.B1(_02264_),
    .Y(_01827_),
    .A1(net283),
    .A2(net676));
 sg13g2_nand2_1 _15537_ (.Y(_02265_),
    .A(\dp.rf.rf[30][8] ),
    .B(net678));
 sg13g2_o21ai_1 _15538_ (.B1(_02265_),
    .Y(_01828_),
    .A1(net280),
    .A2(net678));
 sg13g2_nand2_1 _15539_ (.Y(_02266_),
    .A(\dp.rf.rf[30][9] ),
    .B(net676));
 sg13g2_o21ai_1 _15540_ (.B1(_02266_),
    .Y(_01829_),
    .A1(net272),
    .A2(net676));
 sg13g2_nand2_1 _15541_ (.Y(_02267_),
    .A(\dp.rf.rf[30][10] ),
    .B(net677));
 sg13g2_o21ai_1 _15542_ (.B1(_02267_),
    .Y(_01830_),
    .A1(net269),
    .A2(net677));
 sg13g2_buf_1 input51 (.A(readdata[26]),
    .X(net51));
 sg13g2_nand2_1 _15544_ (.Y(_02269_),
    .A(\dp.rf.rf[30][11] ),
    .B(net677));
 sg13g2_o21ai_1 _15545_ (.B1(_02269_),
    .Y(_01831_),
    .A1(net262),
    .A2(net678));
 sg13g2_nand2_1 _15546_ (.Y(_02270_),
    .A(\dp.rf.rf[30][12] ),
    .B(net675));
 sg13g2_o21ai_1 _15547_ (.B1(_02270_),
    .Y(_01832_),
    .A1(net256),
    .A2(net675));
 sg13g2_mux2_1 _15548_ (.A0(\dp.rf.rf[30][13] ),
    .A1(net252),
    .S(_02260_),
    .X(_01833_));
 sg13g2_buf_1 input50 (.A(readdata[25]),
    .X(net50));
 sg13g2_nand2_1 _15550_ (.Y(_02272_),
    .A(\dp.rf.rf[30][14] ),
    .B(net674));
 sg13g2_o21ai_1 _15551_ (.B1(_02272_),
    .Y(_01834_),
    .A1(net248),
    .A2(net674));
 sg13g2_nand2_1 _15552_ (.Y(_02273_),
    .A(\dp.rf.rf[30][15] ),
    .B(net675));
 sg13g2_o21ai_1 _15553_ (.B1(_02273_),
    .Y(_01835_),
    .A1(net241),
    .A2(net675));
 sg13g2_nand2_1 _15554_ (.Y(_02274_),
    .A(\dp.rf.rf[30][16] ),
    .B(net676));
 sg13g2_o21ai_1 _15555_ (.B1(_02274_),
    .Y(_01836_),
    .A1(net235),
    .A2(net676));
 sg13g2_nand2_1 _15556_ (.Y(_02275_),
    .A(\dp.rf.rf[30][17] ),
    .B(net673));
 sg13g2_o21ai_1 _15557_ (.B1(_02275_),
    .Y(_01837_),
    .A1(net231),
    .A2(net673));
 sg13g2_nand2_1 _15558_ (.Y(_02276_),
    .A(\dp.rf.rf[30][18] ),
    .B(net672));
 sg13g2_o21ai_1 _15559_ (.B1(_02276_),
    .Y(_01838_),
    .A1(net226),
    .A2(net674));
 sg13g2_nand2_1 _15560_ (.Y(_02277_),
    .A(\dp.rf.rf[30][19] ),
    .B(net672));
 sg13g2_o21ai_1 _15561_ (.B1(_02277_),
    .Y(_01839_),
    .A1(net221),
    .A2(net672));
 sg13g2_nand2_1 _15562_ (.Y(_02278_),
    .A(\dp.rf.rf[30][20] ),
    .B(net673));
 sg13g2_o21ai_1 _15563_ (.B1(_02278_),
    .Y(_01840_),
    .A1(net216),
    .A2(net673));
 sg13g2_nand2_1 _15564_ (.Y(_02279_),
    .A(\dp.rf.rf[30][21] ),
    .B(net671));
 sg13g2_o21ai_1 _15565_ (.B1(_02279_),
    .Y(_01841_),
    .A1(net212),
    .A2(net671));
 sg13g2_nor2_1 _15566_ (.A(\dp.rf.rf[30][22] ),
    .B(_02260_),
    .Y(_02280_));
 sg13g2_a21oi_1 _15567_ (.A1(net207),
    .A2(_02260_),
    .Y(_01842_),
    .B1(_02280_));
 sg13g2_nand2_1 _15568_ (.Y(_02281_),
    .A(\dp.rf.rf[30][23] ),
    .B(net671));
 sg13g2_o21ai_1 _15569_ (.B1(_02281_),
    .Y(_01843_),
    .A1(net200),
    .A2(net671));
 sg13g2_nand2_1 _15570_ (.Y(_02282_),
    .A(\dp.rf.rf[30][24] ),
    .B(net673));
 sg13g2_o21ai_1 _15571_ (.B1(_02282_),
    .Y(_01844_),
    .A1(net197),
    .A2(net673));
 sg13g2_nand2_1 _15572_ (.Y(_02283_),
    .A(\dp.rf.rf[30][25] ),
    .B(net670));
 sg13g2_o21ai_1 _15573_ (.B1(_02283_),
    .Y(_01845_),
    .A1(net189),
    .A2(net670));
 sg13g2_nand2_1 _15574_ (.Y(_02284_),
    .A(\dp.rf.rf[30][26] ),
    .B(net670));
 sg13g2_o21ai_1 _15575_ (.B1(_02284_),
    .Y(_01846_),
    .A1(net184),
    .A2(net670));
 sg13g2_nand2_1 _15576_ (.Y(_02285_),
    .A(\dp.rf.rf[30][27] ),
    .B(net670));
 sg13g2_o21ai_1 _15577_ (.B1(_02285_),
    .Y(_01847_),
    .A1(net180),
    .A2(net670));
 sg13g2_nand2_1 _15578_ (.Y(_02286_),
    .A(\dp.rf.rf[30][28] ),
    .B(net670));
 sg13g2_o21ai_1 _15579_ (.B1(_02286_),
    .Y(_01848_),
    .A1(net306),
    .A2(net670));
 sg13g2_nor2_1 _15580_ (.A(\dp.rf.rf[30][29] ),
    .B(_02260_),
    .Y(_02287_));
 sg13g2_a21oi_1 _15581_ (.A1(net174),
    .A2(_02260_),
    .Y(_01849_),
    .B1(_02287_));
 sg13g2_nand2_1 _15582_ (.Y(_02288_),
    .A(\dp.rf.rf[30][30] ),
    .B(net673));
 sg13g2_o21ai_1 _15583_ (.B1(_02288_),
    .Y(_01850_),
    .A1(net173),
    .A2(net673));
 sg13g2_nand2_1 _15584_ (.Y(_02289_),
    .A(\dp.rf.rf[30][31] ),
    .B(net672));
 sg13g2_o21ai_1 _15585_ (.B1(_02289_),
    .Y(_01851_),
    .A1(net166),
    .A2(net672));
 sg13g2_nor2_1 _15586_ (.A(_08016_),
    .B(_08468_),
    .Y(_02290_));
 sg13g2_buf_1 input49 (.A(readdata[24]),
    .X(net49));
 sg13g2_buf_1 input48 (.A(readdata[23]),
    .X(net48));
 sg13g2_nor2_1 _15589_ (.A(\dp.rf.rf[24][0] ),
    .B(_02290_),
    .Y(_02293_));
 sg13g2_a21oi_1 _15590_ (.A1(net302),
    .A2(net669),
    .Y(_01852_),
    .B1(_02293_));
 sg13g2_or2_1 _15591_ (.X(_02294_),
    .B(_08468_),
    .A(_08016_));
 sg13g2_buf_1 input47 (.A(readdata[22]),
    .X(net47));
 sg13g2_buf_1 input46 (.A(readdata[21]),
    .X(net46));
 sg13g2_buf_1 input45 (.A(readdata[20]),
    .X(net45));
 sg13g2_nand2_1 _15595_ (.Y(_02298_),
    .A(\dp.rf.rf[24][1] ),
    .B(net665));
 sg13g2_o21ai_1 _15596_ (.B1(_02298_),
    .Y(_01853_),
    .A1(net298),
    .A2(net665));
 sg13g2_nand2_1 _15597_ (.Y(_02299_),
    .A(\dp.rf.rf[24][2] ),
    .B(net665));
 sg13g2_o21ai_1 _15598_ (.B1(_02299_),
    .Y(_01854_),
    .A1(net322),
    .A2(net666));
 sg13g2_nand2_1 _15599_ (.Y(_02300_),
    .A(\dp.rf.rf[24][3] ),
    .B(net665));
 sg13g2_o21ai_1 _15600_ (.B1(_02300_),
    .Y(_01855_),
    .A1(net318),
    .A2(net665));
 sg13g2_mux2_1 _15601_ (.A0(\dp.rf.rf[24][4] ),
    .A1(net290),
    .S(net669),
    .X(_01856_));
 sg13g2_nand2_1 _15602_ (.Y(_02301_),
    .A(\dp.rf.rf[24][5] ),
    .B(net663));
 sg13g2_o21ai_1 _15603_ (.B1(_02301_),
    .Y(_01857_),
    .A1(net313),
    .A2(net663));
 sg13g2_nand2_1 _15604_ (.Y(_02302_),
    .A(\dp.rf.rf[24][6] ),
    .B(net664));
 sg13g2_o21ai_1 _15605_ (.B1(_02302_),
    .Y(_01858_),
    .A1(net288),
    .A2(net664));
 sg13g2_nand2_1 _15606_ (.Y(_02303_),
    .A(\dp.rf.rf[24][7] ),
    .B(net664));
 sg13g2_o21ai_1 _15607_ (.B1(_02303_),
    .Y(_01859_),
    .A1(net284),
    .A2(net664));
 sg13g2_nand2_1 _15608_ (.Y(_02304_),
    .A(\dp.rf.rf[24][8] ),
    .B(net666));
 sg13g2_o21ai_1 _15609_ (.B1(_02304_),
    .Y(_01860_),
    .A1(net278),
    .A2(net666));
 sg13g2_buf_1 input44 (.A(readdata[1]),
    .X(net44));
 sg13g2_nand2_1 _15611_ (.Y(_02306_),
    .A(\dp.rf.rf[24][9] ),
    .B(net663));
 sg13g2_o21ai_1 _15612_ (.B1(_02306_),
    .Y(_01861_),
    .A1(net271),
    .A2(net663));
 sg13g2_nand2_1 _15613_ (.Y(_02307_),
    .A(\dp.rf.rf[24][10] ),
    .B(net665));
 sg13g2_o21ai_1 _15614_ (.B1(_02307_),
    .Y(_01862_),
    .A1(net268),
    .A2(net665));
 sg13g2_nand2_1 _15615_ (.Y(_02308_),
    .A(\dp.rf.rf[24][11] ),
    .B(net666));
 sg13g2_o21ai_1 _15616_ (.B1(_02308_),
    .Y(_01863_),
    .A1(net265),
    .A2(net665));
 sg13g2_buf_1 input43 (.A(readdata[19]),
    .X(net43));
 sg13g2_nand2_1 _15618_ (.Y(_02310_),
    .A(\dp.rf.rf[24][12] ),
    .B(net664));
 sg13g2_o21ai_1 _15619_ (.B1(_02310_),
    .Y(_01864_),
    .A1(net258),
    .A2(net664));
 sg13g2_mux2_1 _15620_ (.A0(\dp.rf.rf[24][13] ),
    .A1(net251),
    .S(net669),
    .X(_01865_));
 sg13g2_nor2_1 _15621_ (.A(\dp.rf.rf[24][14] ),
    .B(net669),
    .Y(_02311_));
 sg13g2_a21oi_1 _15622_ (.A1(net247),
    .A2(net669),
    .Y(_01866_),
    .B1(_02311_));
 sg13g2_nand2_1 _15623_ (.Y(_02312_),
    .A(\dp.rf.rf[24][15] ),
    .B(net663));
 sg13g2_o21ai_1 _15624_ (.B1(_02312_),
    .Y(_01867_),
    .A1(net240),
    .A2(net663));
 sg13g2_nand2_1 _15625_ (.Y(_02313_),
    .A(\dp.rf.rf[24][16] ),
    .B(net663));
 sg13g2_o21ai_1 _15626_ (.B1(_02313_),
    .Y(_01868_),
    .A1(net235),
    .A2(net663));
 sg13g2_nor2_1 _15627_ (.A(\dp.rf.rf[24][17] ),
    .B(net669),
    .Y(_02314_));
 sg13g2_a21oi_1 _15628_ (.A1(net231),
    .A2(net669),
    .Y(_01869_),
    .B1(_02314_));
 sg13g2_nand2_1 _15629_ (.Y(_02315_),
    .A(\dp.rf.rf[24][18] ),
    .B(net662));
 sg13g2_o21ai_1 _15630_ (.B1(_02315_),
    .Y(_01870_),
    .A1(net226),
    .A2(net662));
 sg13g2_nand2_1 _15631_ (.Y(_02316_),
    .A(\dp.rf.rf[24][19] ),
    .B(net662));
 sg13g2_o21ai_1 _15632_ (.B1(_02316_),
    .Y(_01871_),
    .A1(net220),
    .A2(net662));
 sg13g2_nor2_1 _15633_ (.A(\dp.rf.rf[24][20] ),
    .B(net668),
    .Y(_02317_));
 sg13g2_a21oi_1 _15634_ (.A1(net217),
    .A2(net668),
    .Y(_01872_),
    .B1(_02317_));
 sg13g2_nand2_1 _15635_ (.Y(_02318_),
    .A(\dp.rf.rf[24][21] ),
    .B(net661));
 sg13g2_o21ai_1 _15636_ (.B1(_02318_),
    .Y(_01873_),
    .A1(net211),
    .A2(net661));
 sg13g2_nor2_1 _15637_ (.A(\dp.rf.rf[24][22] ),
    .B(net668),
    .Y(_02319_));
 sg13g2_a21oi_1 _15638_ (.A1(net207),
    .A2(net668),
    .Y(_01874_),
    .B1(_02319_));
 sg13g2_nand2_1 _15639_ (.Y(_02320_),
    .A(\dp.rf.rf[24][23] ),
    .B(net660));
 sg13g2_o21ai_1 _15640_ (.B1(_02320_),
    .Y(_01875_),
    .A1(net201),
    .A2(net660));
 sg13g2_nand2_1 _15641_ (.Y(_02321_),
    .A(\dp.rf.rf[24][24] ),
    .B(net667));
 sg13g2_o21ai_1 _15642_ (.B1(_02321_),
    .Y(_01876_),
    .A1(net197),
    .A2(net667));
 sg13g2_nand2_1 _15643_ (.Y(_02322_),
    .A(\dp.rf.rf[24][25] ),
    .B(net660));
 sg13g2_o21ai_1 _15644_ (.B1(_02322_),
    .Y(_01877_),
    .A1(net190),
    .A2(net660));
 sg13g2_nand2_1 _15645_ (.Y(_02323_),
    .A(\dp.rf.rf[24][26] ),
    .B(net660));
 sg13g2_o21ai_1 _15646_ (.B1(_02323_),
    .Y(_01878_),
    .A1(net183),
    .A2(net660));
 sg13g2_nand2_1 _15647_ (.Y(_02324_),
    .A(\dp.rf.rf[24][27] ),
    .B(net660));
 sg13g2_o21ai_1 _15648_ (.B1(_02324_),
    .Y(_01879_),
    .A1(net180),
    .A2(net660));
 sg13g2_nand2_1 _15649_ (.Y(_02325_),
    .A(\dp.rf.rf[24][28] ),
    .B(net661));
 sg13g2_o21ai_1 _15650_ (.B1(_02325_),
    .Y(_01880_),
    .A1(net308),
    .A2(net661));
 sg13g2_nor2_1 _15651_ (.A(\dp.rf.rf[24][29] ),
    .B(net668),
    .Y(_02326_));
 sg13g2_a21oi_1 _15652_ (.A1(net175),
    .A2(net668),
    .Y(_01881_),
    .B1(_02326_));
 sg13g2_nor2_1 _15653_ (.A(\dp.rf.rf[24][30] ),
    .B(net668),
    .Y(_02327_));
 sg13g2_a21oi_1 _15654_ (.A1(net172),
    .A2(net668),
    .Y(_01882_),
    .B1(_02327_));
 sg13g2_nand2_1 _15655_ (.Y(_02328_),
    .A(\dp.rf.rf[24][31] ),
    .B(net662));
 sg13g2_o21ai_1 _15656_ (.B1(_02328_),
    .Y(_01883_),
    .A1(net166),
    .A2(net662));
 sg13g2_nand2_1 _15657_ (.Y(_02329_),
    .A(_07396_),
    .B(_08191_));
 sg13g2_buf_1 input42 (.A(readdata[18]),
    .X(net42));
 sg13g2_buf_1 input41 (.A(readdata[17]),
    .X(net41));
 sg13g2_buf_1 input40 (.A(readdata[16]),
    .X(net40));
 sg13g2_nand2_1 _15661_ (.Y(_02333_),
    .A(\dp.rf.rf[23][0] ),
    .B(net449));
 sg13g2_o21ai_1 _15662_ (.B1(_02333_),
    .Y(_01884_),
    .A1(net301),
    .A2(net449));
 sg13g2_nand2_1 _15663_ (.Y(_02334_),
    .A(\dp.rf.rf[23][1] ),
    .B(net454));
 sg13g2_o21ai_1 _15664_ (.B1(_02334_),
    .Y(_01885_),
    .A1(net298),
    .A2(net454));
 sg13g2_nand2_1 _15665_ (.Y(_02335_),
    .A(\dp.rf.rf[23][2] ),
    .B(net455));
 sg13g2_o21ai_1 _15666_ (.B1(_02335_),
    .Y(_01886_),
    .A1(net324),
    .A2(net455));
 sg13g2_nand2_1 _15667_ (.Y(_02336_),
    .A(\dp.rf.rf[23][3] ),
    .B(net454));
 sg13g2_o21ai_1 _15668_ (.B1(_02336_),
    .Y(_01887_),
    .A1(net319),
    .A2(net454));
 sg13g2_mux2_1 _15669_ (.A0(net292),
    .A1(\dp.rf.rf[23][4] ),
    .S(net451),
    .X(_01888_));
 sg13g2_nand2_1 _15670_ (.Y(_02337_),
    .A(\dp.rf.rf[23][5] ),
    .B(net453));
 sg13g2_o21ai_1 _15671_ (.B1(_02337_),
    .Y(_01889_),
    .A1(net313),
    .A2(net453));
 sg13g2_nand2_1 _15672_ (.Y(_02338_),
    .A(\dp.rf.rf[23][6] ),
    .B(net453));
 sg13g2_o21ai_1 _15673_ (.B1(_02338_),
    .Y(_01890_),
    .A1(net287),
    .A2(net453));
 sg13g2_nand2_1 _15674_ (.Y(_02339_),
    .A(\dp.rf.rf[23][7] ),
    .B(net452));
 sg13g2_o21ai_1 _15675_ (.B1(_02339_),
    .Y(_01891_),
    .A1(net281),
    .A2(net452));
 sg13g2_nand2_1 _15676_ (.Y(_02340_),
    .A(\dp.rf.rf[23][8] ),
    .B(net455));
 sg13g2_o21ai_1 _15677_ (.B1(_02340_),
    .Y(_01892_),
    .A1(net279),
    .A2(net455));
 sg13g2_buf_1 input39 (.A(readdata[15]),
    .X(net39));
 sg13g2_nand2_1 _15679_ (.Y(_02342_),
    .A(\dp.rf.rf[23][9] ),
    .B(net452));
 sg13g2_o21ai_1 _15680_ (.B1(_02342_),
    .Y(_01893_),
    .A1(net272),
    .A2(net452));
 sg13g2_nand2_1 _15681_ (.Y(_02343_),
    .A(\dp.rf.rf[23][10] ),
    .B(net454));
 sg13g2_o21ai_1 _15682_ (.B1(_02343_),
    .Y(_01894_),
    .A1(net269),
    .A2(net454));
 sg13g2_buf_1 input38 (.A(readdata[14]),
    .X(net38));
 sg13g2_nand2_1 _15684_ (.Y(_02345_),
    .A(\dp.rf.rf[23][11] ),
    .B(net454));
 sg13g2_o21ai_1 _15685_ (.B1(_02345_),
    .Y(_01895_),
    .A1(net264),
    .A2(net454));
 sg13g2_nand2_1 _15686_ (.Y(_02346_),
    .A(\dp.rf.rf[23][12] ),
    .B(net452));
 sg13g2_o21ai_1 _15687_ (.B1(_02346_),
    .Y(_01896_),
    .A1(net256),
    .A2(net452));
 sg13g2_mux2_1 _15688_ (.A0(net253),
    .A1(\dp.rf.rf[23][13] ),
    .S(net455),
    .X(_01897_));
 sg13g2_nand2_1 _15689_ (.Y(_02347_),
    .A(\dp.rf.rf[23][14] ),
    .B(net448));
 sg13g2_o21ai_1 _15690_ (.B1(_02347_),
    .Y(_01898_),
    .A1(net246),
    .A2(net448));
 sg13g2_nand2_1 _15691_ (.Y(_02348_),
    .A(\dp.rf.rf[23][15] ),
    .B(net453));
 sg13g2_o21ai_1 _15692_ (.B1(_02348_),
    .Y(_01899_),
    .A1(net241),
    .A2(net453));
 sg13g2_nand2_1 _15693_ (.Y(_02349_),
    .A(\dp.rf.rf[23][16] ),
    .B(net452));
 sg13g2_o21ai_1 _15694_ (.B1(_02349_),
    .Y(_01900_),
    .A1(net237),
    .A2(net452));
 sg13g2_nand2_1 _15695_ (.Y(_02350_),
    .A(\dp.rf.rf[23][17] ),
    .B(net451));
 sg13g2_o21ai_1 _15696_ (.B1(_02350_),
    .Y(_01901_),
    .A1(net232),
    .A2(net451));
 sg13g2_nand2_1 _15697_ (.Y(_02351_),
    .A(\dp.rf.rf[23][18] ),
    .B(net451));
 sg13g2_o21ai_1 _15698_ (.B1(_02351_),
    .Y(_01902_),
    .A1(net224),
    .A2(net451));
 sg13g2_nand2_1 _15699_ (.Y(_02352_),
    .A(\dp.rf.rf[23][19] ),
    .B(net449));
 sg13g2_o21ai_1 _15700_ (.B1(_02352_),
    .Y(_01903_),
    .A1(net223),
    .A2(net449));
 sg13g2_buf_1 input37 (.A(readdata[13]),
    .X(net37));
 sg13g2_nand2_1 _15702_ (.Y(_02354_),
    .A(\dp.rf.rf[23][20] ),
    .B(net448));
 sg13g2_o21ai_1 _15703_ (.B1(_02354_),
    .Y(_01904_),
    .A1(net216),
    .A2(net448));
 sg13g2_nand2_1 _15704_ (.Y(_02355_),
    .A(\dp.rf.rf[23][21] ),
    .B(net448));
 sg13g2_o21ai_1 _15705_ (.B1(_02355_),
    .Y(_01905_),
    .A1(net212),
    .A2(net448));
 sg13g2_buf_1 input36 (.A(readdata[12]),
    .X(net36));
 sg13g2_nand2_1 _15707_ (.Y(_02357_),
    .A(\dp.rf.rf[23][22] ),
    .B(net450));
 sg13g2_o21ai_1 _15708_ (.B1(_02357_),
    .Y(_01906_),
    .A1(net207),
    .A2(net450));
 sg13g2_nand2_1 _15709_ (.Y(_02358_),
    .A(\dp.rf.rf[23][23] ),
    .B(net447));
 sg13g2_o21ai_1 _15710_ (.B1(_02358_),
    .Y(_01907_),
    .A1(net200),
    .A2(net447));
 sg13g2_nand2_1 _15711_ (.Y(_02359_),
    .A(\dp.rf.rf[23][24] ),
    .B(net450));
 sg13g2_o21ai_1 _15712_ (.B1(_02359_),
    .Y(_01908_),
    .A1(net198),
    .A2(net450));
 sg13g2_nand2_1 _15713_ (.Y(_02360_),
    .A(\dp.rf.rf[23][25] ),
    .B(net447));
 sg13g2_o21ai_1 _15714_ (.B1(_02360_),
    .Y(_01909_),
    .A1(net189),
    .A2(net447));
 sg13g2_nand2_1 _15715_ (.Y(_02361_),
    .A(\dp.rf.rf[23][26] ),
    .B(net447));
 sg13g2_o21ai_1 _15716_ (.B1(_02361_),
    .Y(_01910_),
    .A1(net183),
    .A2(net447));
 sg13g2_nand2_1 _15717_ (.Y(_02362_),
    .A(\dp.rf.rf[23][27] ),
    .B(net447));
 sg13g2_o21ai_1 _15718_ (.B1(_02362_),
    .Y(_01911_),
    .A1(net179),
    .A2(net447));
 sg13g2_nand2_1 _15719_ (.Y(_02363_),
    .A(\dp.rf.rf[23][28] ),
    .B(net448));
 sg13g2_o21ai_1 _15720_ (.B1(_02363_),
    .Y(_01912_),
    .A1(net307),
    .A2(net448));
 sg13g2_nand2_1 _15721_ (.Y(_02364_),
    .A(\dp.rf.rf[23][29] ),
    .B(net450));
 sg13g2_o21ai_1 _15722_ (.B1(_02364_),
    .Y(_01913_),
    .A1(net174),
    .A2(net450));
 sg13g2_nand2_1 _15723_ (.Y(_02365_),
    .A(\dp.rf.rf[23][30] ),
    .B(net450));
 sg13g2_o21ai_1 _15724_ (.B1(_02365_),
    .Y(_01914_),
    .A1(net172),
    .A2(net450));
 sg13g2_nand2_1 _15725_ (.Y(_02366_),
    .A(\dp.rf.rf[23][31] ),
    .B(net449));
 sg13g2_o21ai_1 _15726_ (.B1(_02366_),
    .Y(_01915_),
    .A1(net165),
    .A2(net449));
 sg13g2_or2_1 _15727_ (.X(_02367_),
    .B(_07787_),
    .A(_02173_));
 sg13g2_buf_1 input35 (.A(readdata[11]),
    .X(net35));
 sg13g2_buf_1 input34 (.A(readdata[10]),
    .X(net34));
 sg13g2_buf_1 input33 (.A(readdata[0]),
    .X(net33));
 sg13g2_nand2_1 _15731_ (.Y(_02371_),
    .A(\dp.rf.rf[31][0] ),
    .B(net437));
 sg13g2_o21ai_1 _15732_ (.B1(_02371_),
    .Y(_01916_),
    .A1(net301),
    .A2(net437));
 sg13g2_nand2_1 _15733_ (.Y(_02372_),
    .A(\dp.rf.rf[31][1] ),
    .B(net444));
 sg13g2_o21ai_1 _15734_ (.B1(_02372_),
    .Y(_01917_),
    .A1(net298),
    .A2(net444));
 sg13g2_nand2_1 _15735_ (.Y(_02373_),
    .A(\dp.rf.rf[31][2] ),
    .B(net445));
 sg13g2_o21ai_1 _15736_ (.B1(_02373_),
    .Y(_01918_),
    .A1(net322),
    .A2(net444));
 sg13g2_nand2_1 _15737_ (.Y(_02374_),
    .A(\dp.rf.rf[31][3] ),
    .B(net444));
 sg13g2_o21ai_1 _15738_ (.B1(_02374_),
    .Y(_01919_),
    .A1(net318),
    .A2(net444));
 sg13g2_mux2_1 _15739_ (.A0(net292),
    .A1(\dp.rf.rf[31][4] ),
    .S(net440),
    .X(_01920_));
 sg13g2_nand2_1 _15740_ (.Y(_02375_),
    .A(\dp.rf.rf[31][5] ),
    .B(net443));
 sg13g2_o21ai_1 _15741_ (.B1(_02375_),
    .Y(_01921_),
    .A1(net312),
    .A2(net443));
 sg13g2_nand2_1 _15742_ (.Y(_02376_),
    .A(\dp.rf.rf[31][6] ),
    .B(net443));
 sg13g2_o21ai_1 _15743_ (.B1(_02376_),
    .Y(_01922_),
    .A1(net288),
    .A2(net443));
 sg13g2_nand2_1 _15744_ (.Y(_02377_),
    .A(\dp.rf.rf[31][7] ),
    .B(net442));
 sg13g2_o21ai_1 _15745_ (.B1(_02377_),
    .Y(_01923_),
    .A1(net283),
    .A2(net442));
 sg13g2_nand2_1 _15746_ (.Y(_02378_),
    .A(\dp.rf.rf[31][8] ),
    .B(net445));
 sg13g2_o21ai_1 _15747_ (.B1(_02378_),
    .Y(_01924_),
    .A1(net278),
    .A2(net445));
 sg13g2_buf_1 input32 (.A(instr[9]),
    .X(net32));
 sg13g2_nand2_1 _15749_ (.Y(_02380_),
    .A(\dp.rf.rf[31][9] ),
    .B(net442));
 sg13g2_o21ai_1 _15750_ (.B1(_02380_),
    .Y(_01925_),
    .A1(net273),
    .A2(net442));
 sg13g2_nand2_1 _15751_ (.Y(_02381_),
    .A(\dp.rf.rf[31][10] ),
    .B(net444));
 sg13g2_o21ai_1 _15752_ (.B1(_02381_),
    .Y(_01926_),
    .A1(net269),
    .A2(net444));
 sg13g2_buf_1 input31 (.A(instr[8]),
    .X(net31));
 sg13g2_nand2_1 _15754_ (.Y(_02383_),
    .A(\dp.rf.rf[31][11] ),
    .B(net444));
 sg13g2_o21ai_1 _15755_ (.B1(_02383_),
    .Y(_01927_),
    .A1(net262),
    .A2(net445));
 sg13g2_nand2_1 _15756_ (.Y(_02384_),
    .A(\dp.rf.rf[31][12] ),
    .B(net443));
 sg13g2_o21ai_1 _15757_ (.B1(_02384_),
    .Y(_01928_),
    .A1(net256),
    .A2(net443));
 sg13g2_mux2_1 _15758_ (.A0(net251),
    .A1(\dp.rf.rf[31][13] ),
    .S(net440),
    .X(_01929_));
 sg13g2_nand2_1 _15759_ (.Y(_02385_),
    .A(\dp.rf.rf[31][14] ),
    .B(net440));
 sg13g2_o21ai_1 _15760_ (.B1(_02385_),
    .Y(_01930_),
    .A1(net248),
    .A2(net440));
 sg13g2_nand2_1 _15761_ (.Y(_02386_),
    .A(\dp.rf.rf[31][15] ),
    .B(net442));
 sg13g2_o21ai_1 _15762_ (.B1(_02386_),
    .Y(_01931_),
    .A1(net241),
    .A2(net442));
 sg13g2_nand2_1 _15763_ (.Y(_02387_),
    .A(\dp.rf.rf[31][16] ),
    .B(net442));
 sg13g2_o21ai_1 _15764_ (.B1(_02387_),
    .Y(_01932_),
    .A1(net234),
    .A2(net442));
 sg13g2_nand2_1 _15765_ (.Y(_02388_),
    .A(\dp.rf.rf[31][17] ),
    .B(net438));
 sg13g2_o21ai_1 _15766_ (.B1(_02388_),
    .Y(_01933_),
    .A1(net231),
    .A2(net438));
 sg13g2_nand2_1 _15767_ (.Y(_02389_),
    .A(\dp.rf.rf[31][18] ),
    .B(net441));
 sg13g2_o21ai_1 _15768_ (.B1(_02389_),
    .Y(_01934_),
    .A1(net224),
    .A2(net441));
 sg13g2_nand2_1 _15769_ (.Y(_02390_),
    .A(\dp.rf.rf[31][19] ),
    .B(net437));
 sg13g2_o21ai_1 _15770_ (.B1(_02390_),
    .Y(_01935_),
    .A1(net221),
    .A2(net437));
 sg13g2_buf_1 input30 (.A(instr[7]),
    .X(net30));
 sg13g2_nand2_1 _15772_ (.Y(_02392_),
    .A(\dp.rf.rf[31][20] ),
    .B(net438));
 sg13g2_o21ai_1 _15773_ (.B1(_02392_),
    .Y(_01936_),
    .A1(net216),
    .A2(net438));
 sg13g2_nand2_1 _15774_ (.Y(_02393_),
    .A(\dp.rf.rf[31][21] ),
    .B(net436));
 sg13g2_o21ai_1 _15775_ (.B1(_02393_),
    .Y(_01937_),
    .A1(net212),
    .A2(net436));
 sg13g2_buf_1 input29 (.A(instr[6]),
    .X(net29));
 sg13g2_nand2_1 _15777_ (.Y(_02395_),
    .A(\dp.rf.rf[31][22] ),
    .B(net439));
 sg13g2_o21ai_1 _15778_ (.B1(_02395_),
    .Y(_01938_),
    .A1(net207),
    .A2(net439));
 sg13g2_nand2_1 _15779_ (.Y(_02396_),
    .A(\dp.rf.rf[31][23] ),
    .B(net435));
 sg13g2_o21ai_1 _15780_ (.B1(_02396_),
    .Y(_01939_),
    .A1(net200),
    .A2(net435));
 sg13g2_nand2_1 _15781_ (.Y(_02397_),
    .A(\dp.rf.rf[31][24] ),
    .B(net438));
 sg13g2_o21ai_1 _15782_ (.B1(_02397_),
    .Y(_01940_),
    .A1(net198),
    .A2(net438));
 sg13g2_nand2_1 _15783_ (.Y(_02398_),
    .A(\dp.rf.rf[31][25] ),
    .B(net435));
 sg13g2_o21ai_1 _15784_ (.B1(_02398_),
    .Y(_01941_),
    .A1(net190),
    .A2(net435));
 sg13g2_nand2_1 _15785_ (.Y(_02399_),
    .A(\dp.rf.rf[31][26] ),
    .B(net435));
 sg13g2_o21ai_1 _15786_ (.B1(_02399_),
    .Y(_01942_),
    .A1(net183),
    .A2(net435));
 sg13g2_nand2_1 _15787_ (.Y(_02400_),
    .A(\dp.rf.rf[31][27] ),
    .B(net435));
 sg13g2_o21ai_1 _15788_ (.B1(_02400_),
    .Y(_01943_),
    .A1(net180),
    .A2(net435));
 sg13g2_nand2_1 _15789_ (.Y(_02401_),
    .A(\dp.rf.rf[31][28] ),
    .B(net436));
 sg13g2_o21ai_1 _15790_ (.B1(_02401_),
    .Y(_01944_),
    .A1(net306),
    .A2(net436));
 sg13g2_nand2_1 _15791_ (.Y(_02402_),
    .A(\dp.rf.rf[31][29] ),
    .B(net438));
 sg13g2_o21ai_1 _15792_ (.B1(_02402_),
    .Y(_01945_),
    .A1(net175),
    .A2(net439));
 sg13g2_nand2_1 _15793_ (.Y(_02403_),
    .A(\dp.rf.rf[31][30] ),
    .B(net438));
 sg13g2_o21ai_1 _15794_ (.B1(_02403_),
    .Y(_01946_),
    .A1(net173),
    .A2(net439));
 sg13g2_nand2_1 _15795_ (.Y(_02404_),
    .A(\dp.rf.rf[31][31] ),
    .B(net437));
 sg13g2_o21ai_1 _15796_ (.B1(_02404_),
    .Y(_01947_),
    .A1(net166),
    .A2(net437));
 sg13g2_nor2_1 _15797_ (.A(_07790_),
    .B(_08201_),
    .Y(_02405_));
 sg13g2_buf_1 input28 (.A(instr[5]),
    .X(net28));
 sg13g2_nor2_1 _15799_ (.A(\dp.rf.rf[21][0] ),
    .B(net433),
    .Y(_02407_));
 sg13g2_a21oi_1 _15800_ (.A1(net302),
    .A2(net433),
    .Y(_01948_),
    .B1(_02407_));
 sg13g2_nand2_2 _15801_ (.Y(_02408_),
    .A(_07795_),
    .B(_08191_));
 sg13g2_buf_2 input27 (.A(instr[4]),
    .X(net27));
 sg13g2_buf_1 input26 (.A(instr[3]),
    .X(net26));
 sg13g2_buf_1 input25 (.A(instr[31]),
    .X(net25));
 sg13g2_nand2_1 _15805_ (.Y(_02412_),
    .A(\dp.rf.rf[21][1] ),
    .B(net431));
 sg13g2_o21ai_1 _15806_ (.B1(_02412_),
    .Y(_01949_),
    .A1(net297),
    .A2(net431));
 sg13g2_nand2_1 _15807_ (.Y(_02413_),
    .A(\dp.rf.rf[21][2] ),
    .B(net432));
 sg13g2_o21ai_1 _15808_ (.B1(_02413_),
    .Y(_01950_),
    .A1(net323),
    .A2(net431));
 sg13g2_nand2_1 _15809_ (.Y(_02414_),
    .A(\dp.rf.rf[21][3] ),
    .B(net431));
 sg13g2_o21ai_1 _15810_ (.B1(_02414_),
    .Y(_01951_),
    .A1(net319),
    .A2(net431));
 sg13g2_mux2_1 _15811_ (.A0(\dp.rf.rf[21][4] ),
    .A1(net293),
    .S(net433),
    .X(_01952_));
 sg13g2_nand2_1 _15812_ (.Y(_02415_),
    .A(\dp.rf.rf[21][5] ),
    .B(net429));
 sg13g2_o21ai_1 _15813_ (.B1(_02415_),
    .Y(_01953_),
    .A1(net313),
    .A2(net429));
 sg13g2_nand2_1 _15814_ (.Y(_02416_),
    .A(\dp.rf.rf[21][6] ),
    .B(net429));
 sg13g2_o21ai_1 _15815_ (.B1(_02416_),
    .Y(_01954_),
    .A1(net287),
    .A2(net429));
 sg13g2_buf_1 input24 (.A(instr[30]),
    .X(net24));
 sg13g2_nand2_1 _15817_ (.Y(_02418_),
    .A(\dp.rf.rf[21][7] ),
    .B(net430));
 sg13g2_o21ai_1 _15818_ (.B1(_02418_),
    .Y(_01955_),
    .A1(net283),
    .A2(net430));
 sg13g2_nand2_1 _15819_ (.Y(_02419_),
    .A(\dp.rf.rf[21][8] ),
    .B(net432));
 sg13g2_o21ai_1 _15820_ (.B1(_02419_),
    .Y(_01956_),
    .A1(net277),
    .A2(net432));
 sg13g2_nand2_1 _15821_ (.Y(_02420_),
    .A(\dp.rf.rf[21][9] ),
    .B(net430));
 sg13g2_o21ai_1 _15822_ (.B1(_02420_),
    .Y(_01957_),
    .A1(net272),
    .A2(net430));
 sg13g2_nand2_1 _15823_ (.Y(_02421_),
    .A(\dp.rf.rf[21][10] ),
    .B(net431));
 sg13g2_o21ai_1 _15824_ (.B1(_02421_),
    .Y(_01958_),
    .A1(net269),
    .A2(net431));
 sg13g2_nand2_1 _15825_ (.Y(_02422_),
    .A(\dp.rf.rf[21][11] ),
    .B(net432));
 sg13g2_o21ai_1 _15826_ (.B1(_02422_),
    .Y(_01959_),
    .A1(net264),
    .A2(net431));
 sg13g2_buf_1 input23 (.A(instr[2]),
    .X(net23));
 sg13g2_nand2_1 _15828_ (.Y(_02424_),
    .A(\dp.rf.rf[21][12] ),
    .B(net429));
 sg13g2_o21ai_1 _15829_ (.B1(_02424_),
    .Y(_01960_),
    .A1(net258),
    .A2(net429));
 sg13g2_mux2_1 _15830_ (.A0(\dp.rf.rf[21][13] ),
    .A1(net252),
    .S(net433),
    .X(_01961_));
 sg13g2_nand2_1 _15831_ (.Y(_02425_),
    .A(\dp.rf.rf[21][14] ),
    .B(net428));
 sg13g2_o21ai_1 _15832_ (.B1(_02425_),
    .Y(_01962_),
    .A1(net245),
    .A2(net428));
 sg13g2_nand2_1 _15833_ (.Y(_02426_),
    .A(\dp.rf.rf[21][15] ),
    .B(net429));
 sg13g2_o21ai_1 _15834_ (.B1(_02426_),
    .Y(_01963_),
    .A1(net241),
    .A2(net429));
 sg13g2_nand2_1 _15835_ (.Y(_02427_),
    .A(\dp.rf.rf[21][16] ),
    .B(net430));
 sg13g2_o21ai_1 _15836_ (.B1(_02427_),
    .Y(_01964_),
    .A1(net237),
    .A2(net430));
 sg13g2_nor2_1 _15837_ (.A(\dp.rf.rf[21][17] ),
    .B(net433),
    .Y(_02428_));
 sg13g2_a21oi_1 _15838_ (.A1(net232),
    .A2(net433),
    .Y(_01965_),
    .B1(_02428_));
 sg13g2_nand2_1 _15839_ (.Y(_02429_),
    .A(\dp.rf.rf[21][18] ),
    .B(net427));
 sg13g2_o21ai_1 _15840_ (.B1(_02429_),
    .Y(_01966_),
    .A1(net224),
    .A2(net427));
 sg13g2_buf_1 input22 (.A(instr[29]),
    .X(net22));
 sg13g2_nand2_1 _15842_ (.Y(_02431_),
    .A(\dp.rf.rf[21][19] ),
    .B(net427));
 sg13g2_o21ai_1 _15843_ (.B1(_02431_),
    .Y(_01967_),
    .A1(net221),
    .A2(net427));
 sg13g2_nand2_1 _15844_ (.Y(_02432_),
    .A(\dp.rf.rf[21][20] ),
    .B(net428));
 sg13g2_o21ai_1 _15845_ (.B1(_02432_),
    .Y(_01968_),
    .A1(net216),
    .A2(net428));
 sg13g2_nand2_1 _15846_ (.Y(_02433_),
    .A(\dp.rf.rf[21][21] ),
    .B(net426));
 sg13g2_o21ai_1 _15847_ (.B1(_02433_),
    .Y(_01969_),
    .A1(net212),
    .A2(net426));
 sg13g2_nor2_1 _15848_ (.A(\dp.rf.rf[21][22] ),
    .B(net434),
    .Y(_02434_));
 sg13g2_a21oi_1 _15849_ (.A1(net207),
    .A2(net434),
    .Y(_01970_),
    .B1(_02434_));
 sg13g2_nand2_1 _15850_ (.Y(_02435_),
    .A(\dp.rf.rf[21][23] ),
    .B(net425));
 sg13g2_o21ai_1 _15851_ (.B1(_02435_),
    .Y(_01971_),
    .A1(net201),
    .A2(net425));
 sg13g2_nand2_1 _15852_ (.Y(_02436_),
    .A(\dp.rf.rf[21][24] ),
    .B(net428));
 sg13g2_o21ai_1 _15853_ (.B1(_02436_),
    .Y(_01972_),
    .A1(net198),
    .A2(net428));
 sg13g2_nand2_1 _15854_ (.Y(_02437_),
    .A(\dp.rf.rf[21][25] ),
    .B(net425));
 sg13g2_o21ai_1 _15855_ (.B1(_02437_),
    .Y(_01973_),
    .A1(net189),
    .A2(net425));
 sg13g2_nand2_1 _15856_ (.Y(_02438_),
    .A(\dp.rf.rf[21][26] ),
    .B(net425));
 sg13g2_o21ai_1 _15857_ (.B1(_02438_),
    .Y(_01974_),
    .A1(net184),
    .A2(net425));
 sg13g2_nand2_1 _15858_ (.Y(_02439_),
    .A(\dp.rf.rf[21][27] ),
    .B(net425));
 sg13g2_o21ai_1 _15859_ (.B1(_02439_),
    .Y(_01975_),
    .A1(net179),
    .A2(net425));
 sg13g2_nand2_1 _15860_ (.Y(_02440_),
    .A(\dp.rf.rf[21][28] ),
    .B(net426));
 sg13g2_o21ai_1 _15861_ (.B1(_02440_),
    .Y(_01976_),
    .A1(net307),
    .A2(net426));
 sg13g2_nor2_1 _15862_ (.A(\dp.rf.rf[21][29] ),
    .B(net433),
    .Y(_02441_));
 sg13g2_a21oi_1 _15863_ (.A1(net174),
    .A2(net433),
    .Y(_01977_),
    .B1(_02441_));
 sg13g2_nor2_1 _15864_ (.A(\dp.rf.rf[21][30] ),
    .B(net434),
    .Y(_02442_));
 sg13g2_a21oi_1 _15865_ (.A1(net173),
    .A2(net434),
    .Y(_01978_),
    .B1(_02442_));
 sg13g2_nand2_1 _15866_ (.Y(_02443_),
    .A(\dp.rf.rf[21][31] ),
    .B(net427));
 sg13g2_o21ai_1 _15867_ (.B1(_02443_),
    .Y(_01979_),
    .A1(net165),
    .A2(net427));
 sg13g2_nand2_1 _15868_ (.Y(_02444_),
    .A(_07930_),
    .B(_08311_));
 sg13g2_buf_1 input21 (.A(instr[28]),
    .X(net21));
 sg13g2_buf_1 input20 (.A(instr[27]),
    .X(net20));
 sg13g2_buf_1 input19 (.A(instr[26]),
    .X(net19));
 sg13g2_nand2_1 _15872_ (.Y(_02448_),
    .A(\dp.rf.rf[6][0] ),
    .B(net657));
 sg13g2_o21ai_1 _15873_ (.B1(_02448_),
    .Y(_01980_),
    .A1(net303),
    .A2(net657));
 sg13g2_nand2_1 _15874_ (.Y(_02449_),
    .A(\dp.rf.rf[6][1] ),
    .B(net659));
 sg13g2_o21ai_1 _15875_ (.B1(_02449_),
    .Y(_01981_),
    .A1(net297),
    .A2(net658));
 sg13g2_nand2_1 _15876_ (.Y(_02450_),
    .A(\dp.rf.rf[6][2] ),
    .B(net659));
 sg13g2_o21ai_1 _15877_ (.B1(_02450_),
    .Y(_01982_),
    .A1(net321),
    .A2(net658));
 sg13g2_nand2_1 _15878_ (.Y(_02451_),
    .A(\dp.rf.rf[6][3] ),
    .B(net658));
 sg13g2_o21ai_1 _15879_ (.B1(_02451_),
    .Y(_01983_),
    .A1(net315),
    .A2(net658));
 sg13g2_mux2_1 _15880_ (.A0(net290),
    .A1(\dp.rf.rf[6][4] ),
    .S(net649),
    .X(_01984_));
 sg13g2_nand2_1 _15881_ (.Y(_02452_),
    .A(\dp.rf.rf[6][5] ),
    .B(net655));
 sg13g2_o21ai_1 _15882_ (.B1(_02452_),
    .Y(_01985_),
    .A1(net311),
    .A2(net655));
 sg13g2_nand2_1 _15883_ (.Y(_02453_),
    .A(\dp.rf.rf[6][6] ),
    .B(net655));
 sg13g2_o21ai_1 _15884_ (.B1(_02453_),
    .Y(_01986_),
    .A1(net285),
    .A2(net655));
 sg13g2_nand2_1 _15885_ (.Y(_02454_),
    .A(\dp.rf.rf[6][7] ),
    .B(net655));
 sg13g2_o21ai_1 _15886_ (.B1(_02454_),
    .Y(_01987_),
    .A1(net282),
    .A2(net655));
 sg13g2_nand2_1 _15887_ (.Y(_02455_),
    .A(\dp.rf.rf[6][8] ),
    .B(net656));
 sg13g2_o21ai_1 _15888_ (.B1(_02455_),
    .Y(_01988_),
    .A1(net276),
    .A2(net658));
 sg13g2_buf_1 input18 (.A(instr[25]),
    .X(net18));
 sg13g2_nand2_1 _15890_ (.Y(_02457_),
    .A(\dp.rf.rf[6][9] ),
    .B(net657));
 sg13g2_o21ai_1 _15891_ (.B1(_02457_),
    .Y(_01989_),
    .A1(net275),
    .A2(net657));
 sg13g2_nand2_1 _15892_ (.Y(_02458_),
    .A(\dp.rf.rf[6][10] ),
    .B(net656));
 sg13g2_o21ai_1 _15893_ (.B1(_02458_),
    .Y(_01990_),
    .A1(net267),
    .A2(net656));
 sg13g2_buf_1 input17 (.A(instr[24]),
    .X(net17));
 sg13g2_nand2_1 _15895_ (.Y(_02460_),
    .A(\dp.rf.rf[6][11] ),
    .B(net658));
 sg13g2_o21ai_1 _15896_ (.B1(_02460_),
    .Y(_01991_),
    .A1(net263),
    .A2(net658));
 sg13g2_nand2_1 _15897_ (.Y(_02461_),
    .A(\dp.rf.rf[6][12] ),
    .B(net656));
 sg13g2_o21ai_1 _15898_ (.B1(_02461_),
    .Y(_01992_),
    .A1(net259),
    .A2(net656));
 sg13g2_mux2_1 _15899_ (.A0(net249),
    .A1(\dp.rf.rf[6][13] ),
    .S(net657),
    .X(_01993_));
 sg13g2_nand2_1 _15900_ (.Y(_02462_),
    .A(\dp.rf.rf[6][14] ),
    .B(net650));
 sg13g2_o21ai_1 _15901_ (.B1(_02462_),
    .Y(_01994_),
    .A1(net245),
    .A2(net650));
 sg13g2_nand2_1 _15902_ (.Y(_02463_),
    .A(\dp.rf.rf[6][15] ),
    .B(net656));
 sg13g2_o21ai_1 _15903_ (.B1(_02463_),
    .Y(_01995_),
    .A1(net243),
    .A2(net656));
 sg13g2_nand2_1 _15904_ (.Y(_02464_),
    .A(\dp.rf.rf[6][16] ),
    .B(net655));
 sg13g2_o21ai_1 _15905_ (.B1(_02464_),
    .Y(_01996_),
    .A1(net236),
    .A2(net655));
 sg13g2_nand2_1 _15906_ (.Y(_02465_),
    .A(\dp.rf.rf[6][17] ),
    .B(net653));
 sg13g2_o21ai_1 _15907_ (.B1(_02465_),
    .Y(_01997_),
    .A1(net230),
    .A2(net650));
 sg13g2_nand2_1 _15908_ (.Y(_02466_),
    .A(\dp.rf.rf[6][18] ),
    .B(net657));
 sg13g2_o21ai_1 _15909_ (.B1(_02466_),
    .Y(_01998_),
    .A1(net225),
    .A2(net657));
 sg13g2_nand2_1 _15910_ (.Y(_02467_),
    .A(\dp.rf.rf[6][19] ),
    .B(net649));
 sg13g2_o21ai_1 _15911_ (.B1(_02467_),
    .Y(_01999_),
    .A1(net223),
    .A2(net649));
 sg13g2_buf_1 input16 (.A(instr[23]),
    .X(net16));
 sg13g2_nand2_1 _15913_ (.Y(_02469_),
    .A(\dp.rf.rf[6][20] ),
    .B(net652));
 sg13g2_o21ai_1 _15914_ (.B1(_02469_),
    .Y(_02000_),
    .A1(net214),
    .A2(net652));
 sg13g2_nand2_1 _15915_ (.Y(_02470_),
    .A(\dp.rf.rf[6][21] ),
    .B(net651));
 sg13g2_o21ai_1 _15916_ (.B1(_02470_),
    .Y(_02001_),
    .A1(net210),
    .A2(net651));
 sg13g2_buf_1 input15 (.A(instr[22]),
    .X(net15));
 sg13g2_nand2_1 _15918_ (.Y(_02472_),
    .A(\dp.rf.rf[6][22] ),
    .B(net652));
 sg13g2_o21ai_1 _15919_ (.B1(_02472_),
    .Y(_02002_),
    .A1(net205),
    .A2(net652));
 sg13g2_nand2_1 _15920_ (.Y(_02473_),
    .A(\dp.rf.rf[6][23] ),
    .B(net649));
 sg13g2_o21ai_1 _15921_ (.B1(_02473_),
    .Y(_02003_),
    .A1(net202),
    .A2(net649));
 sg13g2_nand2_1 _15922_ (.Y(_02474_),
    .A(\dp.rf.rf[6][24] ),
    .B(net651));
 sg13g2_o21ai_1 _15923_ (.B1(_02474_),
    .Y(_02004_),
    .A1(net195),
    .A2(net651));
 sg13g2_nand2_1 _15924_ (.Y(_02475_),
    .A(\dp.rf.rf[6][25] ),
    .B(net651));
 sg13g2_o21ai_1 _15925_ (.B1(_02475_),
    .Y(_02005_),
    .A1(net191),
    .A2(net651));
 sg13g2_nand2_1 _15926_ (.Y(_02476_),
    .A(\dp.rf.rf[6][26] ),
    .B(net652));
 sg13g2_o21ai_1 _15927_ (.B1(_02476_),
    .Y(_02006_),
    .A1(net187),
    .A2(net652));
 sg13g2_nand2_1 _15928_ (.Y(_02477_),
    .A(\dp.rf.rf[6][27] ),
    .B(net649));
 sg13g2_o21ai_1 _15929_ (.B1(_02477_),
    .Y(_02007_),
    .A1(net182),
    .A2(net650));
 sg13g2_nand2_1 _15930_ (.Y(_02478_),
    .A(\dp.rf.rf[6][28] ),
    .B(net651));
 sg13g2_o21ai_1 _15931_ (.B1(_02478_),
    .Y(_02008_),
    .A1(net305),
    .A2(net651));
 sg13g2_nand2_1 _15932_ (.Y(_02479_),
    .A(\dp.rf.rf[6][29] ),
    .B(net653));
 sg13g2_o21ai_1 _15933_ (.B1(_02479_),
    .Y(_02009_),
    .A1(net178),
    .A2(net653));
 sg13g2_nand2_1 _15934_ (.Y(_02480_),
    .A(\dp.rf.rf[6][30] ),
    .B(net652));
 sg13g2_o21ai_1 _15935_ (.B1(_02480_),
    .Y(_02010_),
    .A1(net171),
    .A2(net652));
 sg13g2_nand2_1 _15936_ (.Y(_02481_),
    .A(\dp.rf.rf[6][31] ),
    .B(net649));
 sg13g2_o21ai_1 _15937_ (.B1(_02481_),
    .Y(_02011_),
    .A1(net168),
    .A2(net649));
 sg13g2_nand2_1 _15938_ (.Y(_02482_),
    .A(_07795_),
    .B(_08311_));
 sg13g2_buf_1 input14 (.A(instr[21]),
    .X(net14));
 sg13g2_buf_1 input13 (.A(instr[20]),
    .X(net13));
 sg13g2_buf_1 input12 (.A(instr[1]),
    .X(net12));
 sg13g2_nand2_1 _15942_ (.Y(_02486_),
    .A(\dp.rf.rf[5][0] ),
    .B(net421));
 sg13g2_o21ai_1 _15943_ (.B1(_02486_),
    .Y(_02012_),
    .A1(net300),
    .A2(net421));
 sg13g2_nand2_1 _15944_ (.Y(_02487_),
    .A(\dp.rf.rf[5][1] ),
    .B(net422));
 sg13g2_o21ai_1 _15945_ (.B1(_02487_),
    .Y(_02013_),
    .A1(net296),
    .A2(net422));
 sg13g2_nand2_1 _15946_ (.Y(_02488_),
    .A(\dp.rf.rf[5][2] ),
    .B(net422));
 sg13g2_o21ai_1 _15947_ (.B1(_02488_),
    .Y(_02014_),
    .A1(net321),
    .A2(net422));
 sg13g2_nand2_1 _15948_ (.Y(_02489_),
    .A(\dp.rf.rf[5][3] ),
    .B(net423));
 sg13g2_o21ai_1 _15949_ (.B1(_02489_),
    .Y(_02015_),
    .A1(net316),
    .A2(net423));
 sg13g2_mux2_1 _15950_ (.A0(net291),
    .A1(\dp.rf.rf[5][4] ),
    .S(net421),
    .X(_02016_));
 sg13g2_nand2_1 _15951_ (.Y(_02490_),
    .A(\dp.rf.rf[5][5] ),
    .B(net420));
 sg13g2_o21ai_1 _15952_ (.B1(_02490_),
    .Y(_02017_),
    .A1(net311),
    .A2(net419));
 sg13g2_nand2_1 _15953_ (.Y(_02491_),
    .A(\dp.rf.rf[5][6] ),
    .B(net419));
 sg13g2_o21ai_1 _15954_ (.B1(_02491_),
    .Y(_02018_),
    .A1(net285),
    .A2(net419));
 sg13g2_nand2_1 _15955_ (.Y(_02492_),
    .A(\dp.rf.rf[5][7] ),
    .B(net419));
 sg13g2_o21ai_1 _15956_ (.B1(_02492_),
    .Y(_02019_),
    .A1(net283),
    .A2(net419));
 sg13g2_nand2_1 _15957_ (.Y(_02493_),
    .A(\dp.rf.rf[5][8] ),
    .B(net422));
 sg13g2_o21ai_1 _15958_ (.B1(_02493_),
    .Y(_02020_),
    .A1(net279),
    .A2(net422));
 sg13g2_buf_1 input11 (.A(instr[19]),
    .X(net11));
 sg13g2_nand2_1 _15960_ (.Y(_02495_),
    .A(\dp.rf.rf[5][9] ),
    .B(net421));
 sg13g2_o21ai_1 _15961_ (.B1(_02495_),
    .Y(_02021_),
    .A1(net275),
    .A2(net421));
 sg13g2_nand2_1 _15962_ (.Y(_02496_),
    .A(\dp.rf.rf[5][10] ),
    .B(net420));
 sg13g2_o21ai_1 _15963_ (.B1(_02496_),
    .Y(_02022_),
    .A1(net266),
    .A2(net420));
 sg13g2_buf_1 input10 (.A(instr[18]),
    .X(net10));
 sg13g2_nand2_1 _15965_ (.Y(_02498_),
    .A(\dp.rf.rf[5][11] ),
    .B(net423));
 sg13g2_o21ai_1 _15966_ (.B1(_02498_),
    .Y(_02023_),
    .A1(net263),
    .A2(net423));
 sg13g2_nand2_1 _15967_ (.Y(_02499_),
    .A(\dp.rf.rf[5][12] ),
    .B(net422));
 sg13g2_o21ai_1 _15968_ (.B1(_02499_),
    .Y(_02024_),
    .A1(net259),
    .A2(net422));
 sg13g2_mux2_1 _15969_ (.A0(net250),
    .A1(\dp.rf.rf[5][13] ),
    .S(net421),
    .X(_02025_));
 sg13g2_nand2_1 _15970_ (.Y(_02500_),
    .A(\dp.rf.rf[5][14] ),
    .B(net415));
 sg13g2_o21ai_1 _15971_ (.B1(_02500_),
    .Y(_02026_),
    .A1(net245),
    .A2(net415));
 sg13g2_nand2_1 _15972_ (.Y(_02501_),
    .A(\dp.rf.rf[5][15] ),
    .B(net419));
 sg13g2_o21ai_1 _15973_ (.B1(_02501_),
    .Y(_02027_),
    .A1(net243),
    .A2(net419));
 sg13g2_nand2_1 _15974_ (.Y(_02502_),
    .A(\dp.rf.rf[5][16] ),
    .B(net420));
 sg13g2_o21ai_1 _15975_ (.B1(_02502_),
    .Y(_02028_),
    .A1(net236),
    .A2(net419));
 sg13g2_nand2_1 _15976_ (.Y(_02503_),
    .A(\dp.rf.rf[5][17] ),
    .B(net414));
 sg13g2_o21ai_1 _15977_ (.B1(_02503_),
    .Y(_02029_),
    .A1(net230),
    .A2(net414));
 sg13g2_nand2_1 _15978_ (.Y(_02504_),
    .A(\dp.rf.rf[5][18] ),
    .B(net421));
 sg13g2_o21ai_1 _15979_ (.B1(_02504_),
    .Y(_02030_),
    .A1(net225),
    .A2(net421));
 sg13g2_nand2_1 _15980_ (.Y(_02505_),
    .A(\dp.rf.rf[5][19] ),
    .B(net415));
 sg13g2_o21ai_1 _15981_ (.B1(_02505_),
    .Y(_02031_),
    .A1(net223),
    .A2(net415));
 sg13g2_buf_1 input9 (.A(instr[17]),
    .X(net9));
 sg13g2_nand2_1 _15983_ (.Y(_02507_),
    .A(\dp.rf.rf[5][20] ),
    .B(net417));
 sg13g2_o21ai_1 _15984_ (.B1(_02507_),
    .Y(_02032_),
    .A1(net214),
    .A2(net417));
 sg13g2_nand2_1 _15985_ (.Y(_02508_),
    .A(\dp.rf.rf[5][21] ),
    .B(net416));
 sg13g2_o21ai_1 _15986_ (.B1(_02508_),
    .Y(_02033_),
    .A1(net210),
    .A2(net416));
 sg13g2_buf_1 input8 (.A(instr[16]),
    .X(net8));
 sg13g2_nand2_1 _15988_ (.Y(_02510_),
    .A(\dp.rf.rf[5][22] ),
    .B(net418));
 sg13g2_o21ai_1 _15989_ (.B1(_02510_),
    .Y(_02034_),
    .A1(net205),
    .A2(net417));
 sg13g2_nand2_1 _15990_ (.Y(_02511_),
    .A(\dp.rf.rf[5][23] ),
    .B(net414));
 sg13g2_o21ai_1 _15991_ (.B1(_02511_),
    .Y(_02035_),
    .A1(net202),
    .A2(net414));
 sg13g2_nand2_1 _15992_ (.Y(_02512_),
    .A(\dp.rf.rf[5][24] ),
    .B(net416));
 sg13g2_o21ai_1 _15993_ (.B1(_02512_),
    .Y(_02036_),
    .A1(net195),
    .A2(net416));
 sg13g2_nand2_1 _15994_ (.Y(_02513_),
    .A(\dp.rf.rf[5][25] ),
    .B(net416));
 sg13g2_o21ai_1 _15995_ (.B1(_02513_),
    .Y(_02037_),
    .A1(net191),
    .A2(net416));
 sg13g2_nand2_1 _15996_ (.Y(_02514_),
    .A(\dp.rf.rf[5][26] ),
    .B(net417));
 sg13g2_o21ai_1 _15997_ (.B1(_02514_),
    .Y(_02038_),
    .A1(net187),
    .A2(net417));
 sg13g2_nand2_1 _15998_ (.Y(_02515_),
    .A(\dp.rf.rf[5][27] ),
    .B(net414));
 sg13g2_o21ai_1 _15999_ (.B1(_02515_),
    .Y(_02039_),
    .A1(net182),
    .A2(net414));
 sg13g2_nand2_1 _16000_ (.Y(_02516_),
    .A(\dp.rf.rf[5][28] ),
    .B(net416));
 sg13g2_o21ai_1 _16001_ (.B1(_02516_),
    .Y(_02040_),
    .A1(net305),
    .A2(net416));
 sg13g2_nand2_1 _16002_ (.Y(_02517_),
    .A(\dp.rf.rf[5][29] ),
    .B(net417));
 sg13g2_o21ai_1 _16003_ (.B1(_02517_),
    .Y(_02041_),
    .A1(net178),
    .A2(net418));
 sg13g2_nand2_1 _16004_ (.Y(_02518_),
    .A(\dp.rf.rf[5][30] ),
    .B(net417));
 sg13g2_o21ai_1 _16005_ (.B1(_02518_),
    .Y(_02042_),
    .A1(net171),
    .A2(net417));
 sg13g2_nand2_1 _16006_ (.Y(_02519_),
    .A(\dp.rf.rf[5][31] ),
    .B(net414));
 sg13g2_o21ai_1 _16007_ (.B1(_02519_),
    .Y(_02043_),
    .A1(net165),
    .A2(net414));
 sg13g2_mux2_1 _16008_ (.A0(_07408_),
    .A1(net100),
    .S(net335),
    .X(_02044_));
 sg13g2_mux2_1 _16009_ (.A0(_07424_),
    .A1(net111),
    .S(net335),
    .X(_02045_));
 sg13g2_nand2_1 _16010_ (.Y(_02520_),
    .A(_07396_),
    .B(_07840_));
 sg13g2_buf_1 input7 (.A(instr[15]),
    .X(net7));
 sg13g2_buf_1 input6 (.A(instr[14]),
    .X(net6));
 sg13g2_buf_1 input5 (.A(instr[13]),
    .X(net5));
 sg13g2_nand2_1 _16014_ (.Y(_02524_),
    .A(\dp.rf.rf[3][0] ),
    .B(net408));
 sg13g2_o21ai_1 _16015_ (.B1(_02524_),
    .Y(_02046_),
    .A1(net301),
    .A2(net408));
 sg13g2_nand2_1 _16016_ (.Y(_02525_),
    .A(\dp.rf.rf[3][1] ),
    .B(net412));
 sg13g2_o21ai_1 _16017_ (.B1(_02525_),
    .Y(_02047_),
    .A1(net296),
    .A2(net412));
 sg13g2_nand2_1 _16018_ (.Y(_02526_),
    .A(\dp.rf.rf[3][2] ),
    .B(net412));
 sg13g2_o21ai_1 _16019_ (.B1(_02526_),
    .Y(_02048_),
    .A1(net321),
    .A2(net412));
 sg13g2_nand2_1 _16020_ (.Y(_02527_),
    .A(\dp.rf.rf[3][3] ),
    .B(net413));
 sg13g2_o21ai_1 _16021_ (.B1(_02527_),
    .Y(_02049_),
    .A1(net315),
    .A2(net413));
 sg13g2_mux2_1 _16022_ (.A0(net294),
    .A1(\dp.rf.rf[3][4] ),
    .S(net411),
    .X(_02050_));
 sg13g2_nand2_1 _16023_ (.Y(_02528_),
    .A(\dp.rf.rf[3][5] ),
    .B(net409));
 sg13g2_o21ai_1 _16024_ (.B1(_02528_),
    .Y(_02051_),
    .A1(net311),
    .A2(net409));
 sg13g2_nand2_1 _16025_ (.Y(_02529_),
    .A(\dp.rf.rf[3][6] ),
    .B(net409));
 sg13g2_o21ai_1 _16026_ (.B1(_02529_),
    .Y(_02052_),
    .A1(net286),
    .A2(net409));
 sg13g2_nand2_1 _16027_ (.Y(_02530_),
    .A(\dp.rf.rf[3][7] ),
    .B(net410));
 sg13g2_o21ai_1 _16028_ (.B1(_02530_),
    .Y(_02053_),
    .A1(net281),
    .A2(net410));
 sg13g2_nand2_1 _16029_ (.Y(_02531_),
    .A(\dp.rf.rf[3][8] ),
    .B(net411));
 sg13g2_o21ai_1 _16030_ (.B1(_02531_),
    .Y(_02054_),
    .A1(net276),
    .A2(net411));
 sg13g2_buf_1 input4 (.A(instr[12]),
    .X(net4));
 sg13g2_nand2_1 _16032_ (.Y(_02533_),
    .A(\dp.rf.rf[3][9] ),
    .B(net408));
 sg13g2_o21ai_1 _16033_ (.B1(_02533_),
    .Y(_02055_),
    .A1(net274),
    .A2(net408));
 sg13g2_nand2_1 _16034_ (.Y(_02534_),
    .A(\dp.rf.rf[3][10] ),
    .B(net410));
 sg13g2_o21ai_1 _16035_ (.B1(_02534_),
    .Y(_02056_),
    .A1(net270),
    .A2(net410));
 sg13g2_buf_1 input3 (.A(instr[11]),
    .X(net3));
 sg13g2_nand2_1 _16037_ (.Y(_02536_),
    .A(\dp.rf.rf[3][11] ),
    .B(net412));
 sg13g2_o21ai_1 _16038_ (.B1(_02536_),
    .Y(_02057_),
    .A1(net260),
    .A2(net412));
 sg13g2_nand2_1 _16039_ (.Y(_02537_),
    .A(\dp.rf.rf[3][12] ),
    .B(net412));
 sg13g2_o21ai_1 _16040_ (.B1(_02537_),
    .Y(_02058_),
    .A1(net254),
    .A2(net412));
 sg13g2_mux2_1 _16041_ (.A0(net252),
    .A1(\dp.rf.rf[3][13] ),
    .S(net413),
    .X(_02059_));
 sg13g2_nand2_1 _16042_ (.Y(_02538_),
    .A(\dp.rf.rf[3][14] ),
    .B(net404));
 sg13g2_o21ai_1 _16043_ (.B1(_02538_),
    .Y(_02060_),
    .A1(net247),
    .A2(net404));
 sg13g2_nand2_1 _16044_ (.Y(_02539_),
    .A(\dp.rf.rf[3][15] ),
    .B(net409));
 sg13g2_o21ai_1 _16045_ (.B1(_02539_),
    .Y(_02061_),
    .A1(net243),
    .A2(net409));
 sg13g2_nand2_1 _16046_ (.Y(_02540_),
    .A(\dp.rf.rf[3][16] ),
    .B(net409));
 sg13g2_o21ai_1 _16047_ (.B1(_02540_),
    .Y(_02062_),
    .A1(net237),
    .A2(net409));
 sg13g2_nand2_1 _16048_ (.Y(_02541_),
    .A(\dp.rf.rf[3][17] ),
    .B(net407));
 sg13g2_o21ai_1 _16049_ (.B1(_02541_),
    .Y(_02063_),
    .A1(net229),
    .A2(net407));
 sg13g2_nand2_1 _16050_ (.Y(_02542_),
    .A(\dp.rf.rf[3][18] ),
    .B(net408));
 sg13g2_o21ai_1 _16051_ (.B1(_02542_),
    .Y(_02064_),
    .A1(net228),
    .A2(net408));
 sg13g2_nand2_1 _16052_ (.Y(_02543_),
    .A(\dp.rf.rf[3][19] ),
    .B(net408));
 sg13g2_o21ai_1 _16053_ (.B1(_02543_),
    .Y(_02065_),
    .A1(net222),
    .A2(net408));
 sg13g2_buf_1 input2 (.A(instr[10]),
    .X(net2));
 sg13g2_nand2_1 _16055_ (.Y(_02545_),
    .A(\dp.rf.rf[3][20] ),
    .B(net406));
 sg13g2_o21ai_1 _16056_ (.B1(_02545_),
    .Y(_02066_),
    .A1(net215),
    .A2(net406));
 sg13g2_nand2_1 _16057_ (.Y(_02546_),
    .A(\dp.rf.rf[3][21] ),
    .B(net405));
 sg13g2_o21ai_1 _16058_ (.B1(_02546_),
    .Y(_02067_),
    .A1(net213),
    .A2(net405));
 sg13g2_buf_1 input1 (.A(instr[0]),
    .X(net1));
 sg13g2_nand2_1 _16060_ (.Y(_02548_),
    .A(\dp.rf.rf[3][22] ),
    .B(net406));
 sg13g2_o21ai_1 _16061_ (.B1(_02548_),
    .Y(_02068_),
    .A1(net206),
    .A2(net406));
 sg13g2_nand2_1 _16062_ (.Y(_02549_),
    .A(\dp.rf.rf[3][23] ),
    .B(net404));
 sg13g2_o21ai_1 _16063_ (.B1(_02549_),
    .Y(_02069_),
    .A1(net203),
    .A2(net404));
 sg13g2_nand2_1 _16064_ (.Y(_02550_),
    .A(\dp.rf.rf[3][24] ),
    .B(net405));
 sg13g2_o21ai_1 _16065_ (.B1(_02550_),
    .Y(_02070_),
    .A1(net196),
    .A2(net405));
 sg13g2_nand2_1 _16066_ (.Y(_02551_),
    .A(\dp.rf.rf[3][25] ),
    .B(net405));
 sg13g2_o21ai_1 _16067_ (.B1(_02551_),
    .Y(_02071_),
    .A1(net192),
    .A2(net405));
 sg13g2_nand2_1 _16068_ (.Y(_02552_),
    .A(\dp.rf.rf[3][26] ),
    .B(net406));
 sg13g2_o21ai_1 _16069_ (.B1(_02552_),
    .Y(_02072_),
    .A1(net186),
    .A2(net406));
 sg13g2_nand2_1 _16070_ (.Y(_02553_),
    .A(\dp.rf.rf[3][27] ),
    .B(net404));
 sg13g2_o21ai_1 _16071_ (.B1(_02553_),
    .Y(_02073_),
    .A1(net182),
    .A2(net404));
 sg13g2_nand2_1 _16072_ (.Y(_02554_),
    .A(\dp.rf.rf[3][28] ),
    .B(net405));
 sg13g2_o21ai_1 _16073_ (.B1(_02554_),
    .Y(_02074_),
    .A1(net307),
    .A2(net405));
 sg13g2_nand2_1 _16074_ (.Y(_02555_),
    .A(\dp.rf.rf[3][29] ),
    .B(net406));
 sg13g2_o21ai_1 _16075_ (.B1(_02555_),
    .Y(_02075_),
    .A1(net177),
    .A2(net407));
 sg13g2_nand2_1 _16076_ (.Y(_02556_),
    .A(\dp.rf.rf[3][30] ),
    .B(net406));
 sg13g2_o21ai_1 _16077_ (.B1(_02556_),
    .Y(_02076_),
    .A1(net171),
    .A2(net407));
 sg13g2_nand2_1 _16078_ (.Y(_02557_),
    .A(\dp.rf.rf[3][31] ),
    .B(net404));
 sg13g2_o21ai_1 _16079_ (.B1(_02557_),
    .Y(_02077_),
    .A1(net169),
    .A2(net404));
 sg13g2_dfrbp_1 _16080_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_01054_),
    .Q_N(_00019_),
    .Q(\dp.rf.rf[19][0] ));
 sg13g2_dfrbp_1 _16081_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01055_),
    .Q_N(_01009_),
    .Q(\dp.rf.rf[19][1] ));
 sg13g2_dfrbp_1 _16082_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01056_),
    .Q_N(_00977_),
    .Q(\dp.rf.rf[19][2] ));
 sg13g2_dfrbp_1 _16083_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01057_),
    .Q_N(_00945_),
    .Q(\dp.rf.rf[19][3] ));
 sg13g2_dfrbp_1 _16084_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01058_),
    .Q_N(_00913_),
    .Q(\dp.rf.rf[19][4] ));
 sg13g2_dfrbp_1 _16085_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_08518_),
    .D(_01059_),
    .Q_N(_00881_),
    .Q(\dp.rf.rf[19][5] ));
 sg13g2_dfrbp_1 _16086_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01060_),
    .Q_N(_00849_),
    .Q(\dp.rf.rf[19][6] ));
 sg13g2_dfrbp_1 _16087_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01061_),
    .Q_N(_00817_),
    .Q(\dp.rf.rf[19][7] ));
 sg13g2_dfrbp_1 _16088_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01062_),
    .Q_N(_00785_),
    .Q(\dp.rf.rf[19][8] ));
 sg13g2_dfrbp_1 _16089_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01063_),
    .Q_N(_00753_),
    .Q(\dp.rf.rf[19][9] ));
 sg13g2_dfrbp_1 _16090_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01064_),
    .Q_N(_00721_),
    .Q(\dp.rf.rf[19][10] ));
 sg13g2_dfrbp_1 _16091_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01065_),
    .Q_N(_00689_),
    .Q(\dp.rf.rf[19][11] ));
 sg13g2_dfrbp_1 _16092_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_08518_),
    .D(_01066_),
    .Q_N(_00657_),
    .Q(\dp.rf.rf[19][12] ));
 sg13g2_dfrbp_1 _16093_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_08518_),
    .D(_01067_),
    .Q_N(_00625_),
    .Q(\dp.rf.rf[19][13] ));
 sg13g2_dfrbp_1 _16094_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(_08518_),
    .D(_01068_),
    .Q_N(_00593_),
    .Q(\dp.rf.rf[19][14] ));
 sg13g2_dfrbp_1 _16095_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01069_),
    .Q_N(_00561_),
    .Q(\dp.rf.rf[19][15] ));
 sg13g2_dfrbp_1 _16096_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01070_),
    .Q_N(_00529_),
    .Q(\dp.rf.rf[19][16] ));
 sg13g2_dfrbp_1 _16097_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(_08518_),
    .D(_01071_),
    .Q_N(_00497_),
    .Q(\dp.rf.rf[19][17] ));
 sg13g2_dfrbp_1 _16098_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(_01072_),
    .Q_N(_00466_),
    .Q(\dp.rf.rf[19][18] ));
 sg13g2_dfrbp_1 _16099_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_01073_),
    .Q_N(_00434_),
    .Q(\dp.rf.rf[19][19] ));
 sg13g2_dfrbp_1 _16100_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01074_),
    .Q_N(_00403_),
    .Q(\dp.rf.rf[19][20] ));
 sg13g2_dfrbp_1 _16101_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01075_),
    .Q_N(_00371_),
    .Q(\dp.rf.rf[19][21] ));
 sg13g2_dfrbp_1 _16102_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(_08518_),
    .D(_01076_),
    .Q_N(_00339_),
    .Q(\dp.rf.rf[19][22] ));
 sg13g2_dfrbp_1 _16103_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_01077_),
    .Q_N(_00307_),
    .Q(\dp.rf.rf[19][23] ));
 sg13g2_dfrbp_1 _16104_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01078_),
    .Q_N(_00275_),
    .Q(\dp.rf.rf[19][24] ));
 sg13g2_dfrbp_1 _16105_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01079_),
    .Q_N(_00243_),
    .Q(\dp.rf.rf[19][25] ));
 sg13g2_dfrbp_1 _16106_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01080_),
    .Q_N(_00211_),
    .Q(\dp.rf.rf[19][26] ));
 sg13g2_dfrbp_1 _16107_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01081_),
    .Q_N(_00179_),
    .Q(\dp.rf.rf[19][27] ));
 sg13g2_dfrbp_1 _16108_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01082_),
    .Q_N(_00147_),
    .Q(\dp.rf.rf[19][28] ));
 sg13g2_dfrbp_1 _16109_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01083_),
    .Q_N(_00115_),
    .Q(\dp.rf.rf[19][29] ));
 sg13g2_dfrbp_1 _16110_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01084_),
    .Q_N(_00083_),
    .Q(\dp.rf.rf[19][30] ));
 sg13g2_dfrbp_1 _16111_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01085_),
    .Q_N(_00051_),
    .Q(\dp.rf.rf[19][31] ));
 sg13g2_dfrbp_1 _16112_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_08518_),
    .D(_01086_),
    .Q_N(_00011_),
    .Q(\dp.rf.rf[11][0] ));
 sg13g2_dfrbp_1 _16113_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01087_),
    .Q_N(_01001_),
    .Q(\dp.rf.rf[11][1] ));
 sg13g2_dfrbp_1 _16114_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01088_),
    .Q_N(_00969_),
    .Q(\dp.rf.rf[11][2] ));
 sg13g2_dfrbp_1 _16115_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(_08518_),
    .D(_01089_),
    .Q_N(_00937_),
    .Q(\dp.rf.rf[11][3] ));
 sg13g2_dfrbp_1 _16116_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_08518_),
    .D(_01090_),
    .Q_N(_00905_),
    .Q(\dp.rf.rf[11][4] ));
 sg13g2_dfrbp_1 _16117_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_08518_),
    .D(_01091_),
    .Q_N(_00873_),
    .Q(\dp.rf.rf[11][5] ));
 sg13g2_dfrbp_1 _16118_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01092_),
    .Q_N(_00841_),
    .Q(\dp.rf.rf[11][6] ));
 sg13g2_dfrbp_1 _16119_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_01093_),
    .Q_N(_00809_),
    .Q(\dp.rf.rf[11][7] ));
 sg13g2_dfrbp_1 _16120_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_01094_),
    .Q_N(_00777_),
    .Q(\dp.rf.rf[11][8] ));
 sg13g2_dfrbp_1 _16121_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01095_),
    .Q_N(_00745_),
    .Q(\dp.rf.rf[11][9] ));
 sg13g2_dfrbp_1 _16122_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01096_),
    .Q_N(_00713_),
    .Q(\dp.rf.rf[11][10] ));
 sg13g2_dfrbp_1 _16123_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01097_),
    .Q_N(_00681_),
    .Q(\dp.rf.rf[11][11] ));
 sg13g2_dfrbp_1 _16124_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_08518_),
    .D(_01098_),
    .Q_N(_00649_),
    .Q(\dp.rf.rf[11][12] ));
 sg13g2_dfrbp_1 _16125_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_08518_),
    .D(_01099_),
    .Q_N(_00617_),
    .Q(\dp.rf.rf[11][13] ));
 sg13g2_dfrbp_1 _16126_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01100_),
    .Q_N(_00585_),
    .Q(\dp.rf.rf[11][14] ));
 sg13g2_dfrbp_1 _16127_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_01101_),
    .Q_N(_00553_),
    .Q(\dp.rf.rf[11][15] ));
 sg13g2_dfrbp_1 _16128_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_08518_),
    .D(_01102_),
    .Q_N(_00521_),
    .Q(\dp.rf.rf[11][16] ));
 sg13g2_dfrbp_1 _16129_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(_08518_),
    .D(_01103_),
    .Q_N(_00489_),
    .Q(\dp.rf.rf[11][17] ));
 sg13g2_dfrbp_1 _16130_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(_01104_),
    .Q_N(_00458_),
    .Q(\dp.rf.rf[11][18] ));
 sg13g2_dfrbp_1 _16131_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(_01105_),
    .Q_N(_00426_),
    .Q(\dp.rf.rf[11][19] ));
 sg13g2_dfrbp_1 _16132_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(_08518_),
    .D(_01106_),
    .Q_N(_00395_),
    .Q(\dp.rf.rf[11][20] ));
 sg13g2_dfrbp_1 _16133_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01107_),
    .Q_N(_00363_),
    .Q(\dp.rf.rf[11][21] ));
 sg13g2_dfrbp_1 _16134_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01108_),
    .Q_N(_00331_),
    .Q(\dp.rf.rf[11][22] ));
 sg13g2_dfrbp_1 _16135_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01109_),
    .Q_N(_00299_),
    .Q(\dp.rf.rf[11][23] ));
 sg13g2_dfrbp_1 _16136_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(_08518_),
    .D(_01110_),
    .Q_N(_00267_),
    .Q(\dp.rf.rf[11][24] ));
 sg13g2_dfrbp_1 _16137_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01111_),
    .Q_N(_00235_),
    .Q(\dp.rf.rf[11][25] ));
 sg13g2_dfrbp_1 _16138_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01112_),
    .Q_N(_00203_),
    .Q(\dp.rf.rf[11][26] ));
 sg13g2_dfrbp_1 _16139_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_01113_),
    .Q_N(_00171_),
    .Q(\dp.rf.rf[11][27] ));
 sg13g2_dfrbp_1 _16140_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01114_),
    .Q_N(_00139_),
    .Q(\dp.rf.rf[11][28] ));
 sg13g2_dfrbp_1 _16141_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01115_),
    .Q_N(_00107_),
    .Q(\dp.rf.rf[11][29] ));
 sg13g2_dfrbp_1 _16142_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01116_),
    .Q_N(_00075_),
    .Q(\dp.rf.rf[11][30] ));
 sg13g2_dfrbp_1 _16143_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_08518_),
    .D(_01117_),
    .Q_N(_00043_),
    .Q(\dp.rf.rf[11][31] ));
 sg13g2_dfrbp_1 _16144_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_01118_),
    .Q_N(_00029_),
    .Q(\dp.rf.rf[29][0] ));
 sg13g2_dfrbp_1 _16145_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01119_),
    .Q_N(_01019_),
    .Q(\dp.rf.rf[29][1] ));
 sg13g2_dfrbp_1 _16146_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01120_),
    .Q_N(_00987_),
    .Q(\dp.rf.rf[29][2] ));
 sg13g2_dfrbp_1 _16147_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(_08518_),
    .D(_01121_),
    .Q_N(_00955_),
    .Q(\dp.rf.rf[29][3] ));
 sg13g2_dfrbp_1 _16148_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01122_),
    .Q_N(_00923_),
    .Q(\dp.rf.rf[29][4] ));
 sg13g2_dfrbp_1 _16149_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01123_),
    .Q_N(_00891_),
    .Q(\dp.rf.rf[29][5] ));
 sg13g2_dfrbp_1 _16150_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01124_),
    .Q_N(_00859_),
    .Q(\dp.rf.rf[29][6] ));
 sg13g2_dfrbp_1 _16151_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01125_),
    .Q_N(_00827_),
    .Q(\dp.rf.rf[29][7] ));
 sg13g2_dfrbp_1 _16152_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01126_),
    .Q_N(_00795_),
    .Q(\dp.rf.rf[29][8] ));
 sg13g2_dfrbp_1 _16153_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_08518_),
    .D(_01127_),
    .Q_N(_00763_),
    .Q(\dp.rf.rf[29][9] ));
 sg13g2_dfrbp_1 _16154_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_08518_),
    .D(_01128_),
    .Q_N(_00731_),
    .Q(\dp.rf.rf[29][10] ));
 sg13g2_dfrbp_1 _16155_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01129_),
    .Q_N(_00699_),
    .Q(\dp.rf.rf[29][11] ));
 sg13g2_dfrbp_1 _16156_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_08518_),
    .D(_01130_),
    .Q_N(_00667_),
    .Q(\dp.rf.rf[29][12] ));
 sg13g2_dfrbp_1 _16157_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(_08518_),
    .D(_01131_),
    .Q_N(_00635_),
    .Q(\dp.rf.rf[29][13] ));
 sg13g2_dfrbp_1 _16158_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(_01132_),
    .Q_N(_00603_),
    .Q(\dp.rf.rf[29][14] ));
 sg13g2_dfrbp_1 _16159_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_08518_),
    .D(_01133_),
    .Q_N(_00571_),
    .Q(\dp.rf.rf[29][15] ));
 sg13g2_dfrbp_1 _16160_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01134_),
    .Q_N(_00539_),
    .Q(\dp.rf.rf[29][16] ));
 sg13g2_dfrbp_1 _16161_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(_08518_),
    .D(_01135_),
    .Q_N(_00507_),
    .Q(\dp.rf.rf[29][17] ));
 sg13g2_dfrbp_1 _16162_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01136_),
    .Q_N(_00476_),
    .Q(\dp.rf.rf[29][18] ));
 sg13g2_dfrbp_1 _16163_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_08518_),
    .D(_01137_),
    .Q_N(_00444_),
    .Q(\dp.rf.rf[29][19] ));
 sg13g2_dfrbp_1 _16164_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(_08518_),
    .D(_01138_),
    .Q_N(_00413_),
    .Q(\dp.rf.rf[29][20] ));
 sg13g2_dfrbp_1 _16165_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01139_),
    .Q_N(_00381_),
    .Q(\dp.rf.rf[29][21] ));
 sg13g2_dfrbp_1 _16166_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01140_),
    .Q_N(_00349_),
    .Q(\dp.rf.rf[29][22] ));
 sg13g2_dfrbp_1 _16167_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01141_),
    .Q_N(_00317_),
    .Q(\dp.rf.rf[29][23] ));
 sg13g2_dfrbp_1 _16168_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(_08518_),
    .D(_01142_),
    .Q_N(_00285_),
    .Q(\dp.rf.rf[29][24] ));
 sg13g2_dfrbp_1 _16169_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01143_),
    .Q_N(_00253_),
    .Q(\dp.rf.rf[29][25] ));
 sg13g2_dfrbp_1 _16170_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(_08518_),
    .D(_01144_),
    .Q_N(_00221_),
    .Q(\dp.rf.rf[29][26] ));
 sg13g2_dfrbp_1 _16171_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(_08518_),
    .D(_01145_),
    .Q_N(_00189_),
    .Q(\dp.rf.rf[29][27] ));
 sg13g2_dfrbp_1 _16172_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_01146_),
    .Q_N(_00157_),
    .Q(\dp.rf.rf[29][28] ));
 sg13g2_dfrbp_1 _16173_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01147_),
    .Q_N(_00125_),
    .Q(\dp.rf.rf[29][29] ));
 sg13g2_dfrbp_1 _16174_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(_08518_),
    .D(_01148_),
    .Q_N(_00093_),
    .Q(\dp.rf.rf[29][30] ));
 sg13g2_dfrbp_1 _16175_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01149_),
    .Q_N(_00061_),
    .Q(\dp.rf.rf[29][31] ));
 sg13g2_dfrbp_1 _16176_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_08518_),
    .D(_01150_),
    .Q_N(_00012_),
    .Q(\dp.rf.rf[12][0] ));
 sg13g2_dfrbp_1 _16177_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_08518_),
    .D(_01151_),
    .Q_N(_01002_),
    .Q(\dp.rf.rf[12][1] ));
 sg13g2_dfrbp_1 _16178_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01152_),
    .Q_N(_00970_),
    .Q(\dp.rf.rf[12][2] ));
 sg13g2_dfrbp_1 _16179_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(_08518_),
    .D(_01153_),
    .Q_N(_00938_),
    .Q(\dp.rf.rf[12][3] ));
 sg13g2_dfrbp_1 _16180_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(_01154_),
    .Q_N(_00906_),
    .Q(\dp.rf.rf[12][4] ));
 sg13g2_dfrbp_1 _16181_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_08518_),
    .D(_01155_),
    .Q_N(_00874_),
    .Q(\dp.rf.rf[12][5] ));
 sg13g2_dfrbp_1 _16182_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_08518_),
    .D(_01156_),
    .Q_N(_00842_),
    .Q(\dp.rf.rf[12][6] ));
 sg13g2_dfrbp_1 _16183_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_08518_),
    .D(_01157_),
    .Q_N(_00810_),
    .Q(\dp.rf.rf[12][7] ));
 sg13g2_dfrbp_1 _16184_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01158_),
    .Q_N(_00778_),
    .Q(\dp.rf.rf[12][8] ));
 sg13g2_dfrbp_1 _16185_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(_01159_),
    .Q_N(_00746_),
    .Q(\dp.rf.rf[12][9] ));
 sg13g2_dfrbp_1 _16186_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01160_),
    .Q_N(_00714_),
    .Q(\dp.rf.rf[12][10] ));
 sg13g2_dfrbp_1 _16187_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01161_),
    .Q_N(_00682_),
    .Q(\dp.rf.rf[12][11] ));
 sg13g2_dfrbp_1 _16188_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01162_),
    .Q_N(_00650_),
    .Q(\dp.rf.rf[12][12] ));
 sg13g2_dfrbp_1 _16189_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_08518_),
    .D(_01163_),
    .Q_N(_00618_),
    .Q(\dp.rf.rf[12][13] ));
 sg13g2_dfrbp_1 _16190_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(_08518_),
    .D(_01164_),
    .Q_N(_00586_),
    .Q(\dp.rf.rf[12][14] ));
 sg13g2_dfrbp_1 _16191_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_08518_),
    .D(_01165_),
    .Q_N(_00554_),
    .Q(\dp.rf.rf[12][15] ));
 sg13g2_dfrbp_1 _16192_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_08518_),
    .D(_01166_),
    .Q_N(_00522_),
    .Q(\dp.rf.rf[12][16] ));
 sg13g2_dfrbp_1 _16193_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(_08518_),
    .D(_01167_),
    .Q_N(_00490_),
    .Q(\dp.rf.rf[12][17] ));
 sg13g2_dfrbp_1 _16194_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01168_),
    .Q_N(_00459_),
    .Q(\dp.rf.rf[12][18] ));
 sg13g2_dfrbp_1 _16195_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_01169_),
    .Q_N(_00427_),
    .Q(\dp.rf.rf[12][19] ));
 sg13g2_dfrbp_1 _16196_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01170_),
    .Q_N(_00396_),
    .Q(\dp.rf.rf[12][20] ));
 sg13g2_dfrbp_1 _16197_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01171_),
    .Q_N(_00364_),
    .Q(\dp.rf.rf[12][21] ));
 sg13g2_dfrbp_1 _16198_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(_08518_),
    .D(_01172_),
    .Q_N(_00332_),
    .Q(\dp.rf.rf[12][22] ));
 sg13g2_dfrbp_1 _16199_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_08518_),
    .D(_01173_),
    .Q_N(_00300_),
    .Q(\dp.rf.rf[12][23] ));
 sg13g2_dfrbp_1 _16200_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01174_),
    .Q_N(_00268_),
    .Q(\dp.rf.rf[12][24] ));
 sg13g2_dfrbp_1 _16201_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01175_),
    .Q_N(_00236_),
    .Q(\dp.rf.rf[12][25] ));
 sg13g2_dfrbp_1 _16202_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01176_),
    .Q_N(_00204_),
    .Q(\dp.rf.rf[12][26] ));
 sg13g2_dfrbp_1 _16203_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01177_),
    .Q_N(_00172_),
    .Q(\dp.rf.rf[12][27] ));
 sg13g2_dfrbp_1 _16204_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01178_),
    .Q_N(_00140_),
    .Q(\dp.rf.rf[12][28] ));
 sg13g2_dfrbp_1 _16205_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01179_),
    .Q_N(_00108_),
    .Q(\dp.rf.rf[12][29] ));
 sg13g2_dfrbp_1 _16206_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01180_),
    .Q_N(_00076_),
    .Q(\dp.rf.rf[12][30] ));
 sg13g2_dfrbp_1 _16207_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01181_),
    .Q_N(_00044_),
    .Q(\dp.rf.rf[12][31] ));
 sg13g2_dfrbp_1 _16208_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_08518_),
    .D(_01182_),
    .Q_N(_00013_),
    .Q(\dp.rf.rf[13][0] ));
 sg13g2_dfrbp_1 _16209_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_08518_),
    .D(_01183_),
    .Q_N(_01003_),
    .Q(\dp.rf.rf[13][1] ));
 sg13g2_dfrbp_1 _16210_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01184_),
    .Q_N(_00971_),
    .Q(\dp.rf.rf[13][2] ));
 sg13g2_dfrbp_1 _16211_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(_08518_),
    .D(_01185_),
    .Q_N(_00939_),
    .Q(\dp.rf.rf[13][3] ));
 sg13g2_dfrbp_1 _16212_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(_01186_),
    .Q_N(_00907_),
    .Q(\dp.rf.rf[13][4] ));
 sg13g2_dfrbp_1 _16213_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_08518_),
    .D(_01187_),
    .Q_N(_00875_),
    .Q(\dp.rf.rf[13][5] ));
 sg13g2_dfrbp_1 _16214_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_08518_),
    .D(_01188_),
    .Q_N(_00843_),
    .Q(\dp.rf.rf[13][6] ));
 sg13g2_dfrbp_1 _16215_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_08518_),
    .D(_01189_),
    .Q_N(_00811_),
    .Q(\dp.rf.rf[13][7] ));
 sg13g2_dfrbp_1 _16216_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_08518_),
    .D(_01190_),
    .Q_N(_00779_),
    .Q(\dp.rf.rf[13][8] ));
 sg13g2_dfrbp_1 _16217_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01191_),
    .Q_N(_00747_),
    .Q(\dp.rf.rf[13][9] ));
 sg13g2_dfrbp_1 _16218_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01192_),
    .Q_N(_00715_),
    .Q(\dp.rf.rf[13][10] ));
 sg13g2_dfrbp_1 _16219_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01193_),
    .Q_N(_00683_),
    .Q(\dp.rf.rf[13][11] ));
 sg13g2_dfrbp_1 _16220_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_08518_),
    .D(_01194_),
    .Q_N(_00651_),
    .Q(\dp.rf.rf[13][12] ));
 sg13g2_dfrbp_1 _16221_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_08518_),
    .D(_01195_),
    .Q_N(_00619_),
    .Q(\dp.rf.rf[13][13] ));
 sg13g2_dfrbp_1 _16222_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(_08518_),
    .D(_01196_),
    .Q_N(_00587_),
    .Q(\dp.rf.rf[13][14] ));
 sg13g2_dfrbp_1 _16223_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_08518_),
    .D(_01197_),
    .Q_N(_00555_),
    .Q(\dp.rf.rf[13][15] ));
 sg13g2_dfrbp_1 _16224_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_08518_),
    .D(_01198_),
    .Q_N(_00523_),
    .Q(\dp.rf.rf[13][16] ));
 sg13g2_dfrbp_1 _16225_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01199_),
    .Q_N(_00491_),
    .Q(\dp.rf.rf[13][17] ));
 sg13g2_dfrbp_1 _16226_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01200_),
    .Q_N(_00460_),
    .Q(\dp.rf.rf[13][18] ));
 sg13g2_dfrbp_1 _16227_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_01201_),
    .Q_N(_00428_),
    .Q(\dp.rf.rf[13][19] ));
 sg13g2_dfrbp_1 _16228_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01202_),
    .Q_N(_00397_),
    .Q(\dp.rf.rf[13][20] ));
 sg13g2_dfrbp_1 _16229_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01203_),
    .Q_N(_00365_),
    .Q(\dp.rf.rf[13][21] ));
 sg13g2_dfrbp_1 _16230_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(_08518_),
    .D(_01204_),
    .Q_N(_00333_),
    .Q(\dp.rf.rf[13][22] ));
 sg13g2_dfrbp_1 _16231_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01205_),
    .Q_N(_00301_),
    .Q(\dp.rf.rf[13][23] ));
 sg13g2_dfrbp_1 _16232_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01206_),
    .Q_N(_00269_),
    .Q(\dp.rf.rf[13][24] ));
 sg13g2_dfrbp_1 _16233_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01207_),
    .Q_N(_00237_),
    .Q(\dp.rf.rf[13][25] ));
 sg13g2_dfrbp_1 _16234_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01208_),
    .Q_N(_00205_),
    .Q(\dp.rf.rf[13][26] ));
 sg13g2_dfrbp_1 _16235_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01209_),
    .Q_N(_00173_),
    .Q(\dp.rf.rf[13][27] ));
 sg13g2_dfrbp_1 _16236_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01210_),
    .Q_N(_00141_),
    .Q(\dp.rf.rf[13][28] ));
 sg13g2_dfrbp_1 _16237_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01211_),
    .Q_N(_00109_),
    .Q(\dp.rf.rf[13][29] ));
 sg13g2_dfrbp_1 _16238_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01212_),
    .Q_N(_00077_),
    .Q(\dp.rf.rf[13][30] ));
 sg13g2_dfrbp_1 _16239_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01213_),
    .Q_N(_00045_),
    .Q(\dp.rf.rf[13][31] ));
 sg13g2_dfrbp_1 _16240_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_08518_),
    .D(_01214_),
    .Q_N(_00014_),
    .Q(\dp.rf.rf[14][0] ));
 sg13g2_dfrbp_1 _16241_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_08518_),
    .D(_01215_),
    .Q_N(_01004_),
    .Q(\dp.rf.rf[14][1] ));
 sg13g2_dfrbp_1 _16242_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01216_),
    .Q_N(_00972_),
    .Q(\dp.rf.rf[14][2] ));
 sg13g2_dfrbp_1 _16243_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(_08518_),
    .D(_01217_),
    .Q_N(_00940_),
    .Q(\dp.rf.rf[14][3] ));
 sg13g2_dfrbp_1 _16244_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_08518_),
    .D(_01218_),
    .Q_N(_00908_),
    .Q(\dp.rf.rf[14][4] ));
 sg13g2_dfrbp_1 _16245_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_08518_),
    .D(_01219_),
    .Q_N(_00876_),
    .Q(\dp.rf.rf[14][5] ));
 sg13g2_dfrbp_1 _16246_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_08518_),
    .D(_01220_),
    .Q_N(_00844_),
    .Q(\dp.rf.rf[14][6] ));
 sg13g2_dfrbp_1 _16247_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_08518_),
    .D(_01221_),
    .Q_N(_00812_),
    .Q(\dp.rf.rf[14][7] ));
 sg13g2_dfrbp_1 _16248_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_01222_),
    .Q_N(_00780_),
    .Q(\dp.rf.rf[14][8] ));
 sg13g2_dfrbp_1 _16249_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01223_),
    .Q_N(_00748_),
    .Q(\dp.rf.rf[14][9] ));
 sg13g2_dfrbp_1 _16250_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01224_),
    .Q_N(_00716_),
    .Q(\dp.rf.rf[14][10] ));
 sg13g2_dfrbp_1 _16251_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01225_),
    .Q_N(_00684_),
    .Q(\dp.rf.rf[14][11] ));
 sg13g2_dfrbp_1 _16252_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01226_),
    .Q_N(_00652_),
    .Q(\dp.rf.rf[14][12] ));
 sg13g2_dfrbp_1 _16253_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_08518_),
    .D(_01227_),
    .Q_N(_00620_),
    .Q(\dp.rf.rf[14][13] ));
 sg13g2_dfrbp_1 _16254_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(_08518_),
    .D(_01228_),
    .Q_N(_00588_),
    .Q(\dp.rf.rf[14][14] ));
 sg13g2_dfrbp_1 _16255_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_08518_),
    .D(_01229_),
    .Q_N(_00556_),
    .Q(\dp.rf.rf[14][15] ));
 sg13g2_dfrbp_1 _16256_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_08518_),
    .D(_01230_),
    .Q_N(_00524_),
    .Q(\dp.rf.rf[14][16] ));
 sg13g2_dfrbp_1 _16257_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01231_),
    .Q_N(_00492_),
    .Q(\dp.rf.rf[14][17] ));
 sg13g2_dfrbp_1 _16258_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01232_),
    .Q_N(_00461_),
    .Q(\dp.rf.rf[14][18] ));
 sg13g2_dfrbp_1 _16259_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_01233_),
    .Q_N(_00429_),
    .Q(\dp.rf.rf[14][19] ));
 sg13g2_dfrbp_1 _16260_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(_08518_),
    .D(_01234_),
    .Q_N(_00398_),
    .Q(\dp.rf.rf[14][20] ));
 sg13g2_dfrbp_1 _16261_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01235_),
    .Q_N(_00366_),
    .Q(\dp.rf.rf[14][21] ));
 sg13g2_dfrbp_1 _16262_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(_08518_),
    .D(_01236_),
    .Q_N(_00334_),
    .Q(\dp.rf.rf[14][22] ));
 sg13g2_dfrbp_1 _16263_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_08518_),
    .D(_01237_),
    .Q_N(_00302_),
    .Q(\dp.rf.rf[14][23] ));
 sg13g2_dfrbp_1 _16264_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01238_),
    .Q_N(_00270_),
    .Q(\dp.rf.rf[14][24] ));
 sg13g2_dfrbp_1 _16265_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01239_),
    .Q_N(_00238_),
    .Q(\dp.rf.rf[14][25] ));
 sg13g2_dfrbp_1 _16266_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01240_),
    .Q_N(_00206_),
    .Q(\dp.rf.rf[14][26] ));
 sg13g2_dfrbp_1 _16267_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01241_),
    .Q_N(_00174_),
    .Q(\dp.rf.rf[14][27] ));
 sg13g2_dfrbp_1 _16268_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01242_),
    .Q_N(_00142_),
    .Q(\dp.rf.rf[14][28] ));
 sg13g2_dfrbp_1 _16269_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01243_),
    .Q_N(_00110_),
    .Q(\dp.rf.rf[14][29] ));
 sg13g2_dfrbp_1 _16270_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01244_),
    .Q_N(_00078_),
    .Q(\dp.rf.rf[14][30] ));
 sg13g2_dfrbp_1 _16271_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_01245_),
    .Q_N(_00046_),
    .Q(\dp.rf.rf[14][31] ));
 sg13g2_dfrbp_1 _16272_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_08518_),
    .D(_01246_),
    .Q_N(_00015_),
    .Q(\dp.rf.rf[15][0] ));
 sg13g2_dfrbp_1 _16273_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_08518_),
    .D(_01247_),
    .Q_N(_01005_),
    .Q(\dp.rf.rf[15][1] ));
 sg13g2_dfrbp_1 _16274_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01248_),
    .Q_N(_00973_),
    .Q(\dp.rf.rf[15][2] ));
 sg13g2_dfrbp_1 _16275_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_01249_),
    .Q_N(_00941_),
    .Q(\dp.rf.rf[15][3] ));
 sg13g2_dfrbp_1 _16276_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_08518_),
    .D(_01250_),
    .Q_N(_00909_),
    .Q(\dp.rf.rf[15][4] ));
 sg13g2_dfrbp_1 _16277_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_08518_),
    .D(_01251_),
    .Q_N(_00877_),
    .Q(\dp.rf.rf[15][5] ));
 sg13g2_dfrbp_1 _16278_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_08518_),
    .D(_01252_),
    .Q_N(_00845_),
    .Q(\dp.rf.rf[15][6] ));
 sg13g2_dfrbp_1 _16279_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_08518_),
    .D(_01253_),
    .Q_N(_00813_),
    .Q(\dp.rf.rf[15][7] ));
 sg13g2_dfrbp_1 _16280_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_08518_),
    .D(_01254_),
    .Q_N(_00781_),
    .Q(\dp.rf.rf[15][8] ));
 sg13g2_dfrbp_1 _16281_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01255_),
    .Q_N(_00749_),
    .Q(\dp.rf.rf[15][9] ));
 sg13g2_dfrbp_1 _16282_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01256_),
    .Q_N(_00717_),
    .Q(\dp.rf.rf[15][10] ));
 sg13g2_dfrbp_1 _16283_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01257_),
    .Q_N(_00685_),
    .Q(\dp.rf.rf[15][11] ));
 sg13g2_dfrbp_1 _16284_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_08518_),
    .D(_01258_),
    .Q_N(_00653_),
    .Q(\dp.rf.rf[15][12] ));
 sg13g2_dfrbp_1 _16285_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_08518_),
    .D(_01259_),
    .Q_N(_00621_),
    .Q(\dp.rf.rf[15][13] ));
 sg13g2_dfrbp_1 _16286_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(_08518_),
    .D(_01260_),
    .Q_N(_00589_),
    .Q(\dp.rf.rf[15][14] ));
 sg13g2_dfrbp_1 _16287_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_08518_),
    .D(_01261_),
    .Q_N(_00557_),
    .Q(\dp.rf.rf[15][15] ));
 sg13g2_dfrbp_1 _16288_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_08518_),
    .D(_01262_),
    .Q_N(_00525_),
    .Q(\dp.rf.rf[15][16] ));
 sg13g2_dfrbp_1 _16289_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01263_),
    .Q_N(_00493_),
    .Q(\dp.rf.rf[15][17] ));
 sg13g2_dfrbp_1 _16290_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(_01264_),
    .Q_N(_00462_),
    .Q(\dp.rf.rf[15][18] ));
 sg13g2_dfrbp_1 _16291_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_01265_),
    .Q_N(_00430_),
    .Q(\dp.rf.rf[15][19] ));
 sg13g2_dfrbp_1 _16292_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01266_),
    .Q_N(_00399_),
    .Q(\dp.rf.rf[15][20] ));
 sg13g2_dfrbp_1 _16293_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01267_),
    .Q_N(_00367_),
    .Q(\dp.rf.rf[15][21] ));
 sg13g2_dfrbp_1 _16294_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(_08518_),
    .D(_01268_),
    .Q_N(_00335_),
    .Q(\dp.rf.rf[15][22] ));
 sg13g2_dfrbp_1 _16295_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_08518_),
    .D(_01269_),
    .Q_N(_00303_),
    .Q(\dp.rf.rf[15][23] ));
 sg13g2_dfrbp_1 _16296_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01270_),
    .Q_N(_00271_),
    .Q(\dp.rf.rf[15][24] ));
 sg13g2_dfrbp_1 _16297_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01271_),
    .Q_N(_00239_),
    .Q(\dp.rf.rf[15][25] ));
 sg13g2_dfrbp_1 _16298_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01272_),
    .Q_N(_00207_),
    .Q(\dp.rf.rf[15][26] ));
 sg13g2_dfrbp_1 _16299_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01273_),
    .Q_N(_00175_),
    .Q(\dp.rf.rf[15][27] ));
 sg13g2_dfrbp_1 _16300_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01274_),
    .Q_N(_00143_),
    .Q(\dp.rf.rf[15][28] ));
 sg13g2_dfrbp_1 _16301_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01275_),
    .Q_N(_00111_),
    .Q(\dp.rf.rf[15][29] ));
 sg13g2_dfrbp_1 _16302_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01276_),
    .Q_N(_00079_),
    .Q(\dp.rf.rf[15][30] ));
 sg13g2_dfrbp_1 _16303_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_01277_),
    .Q_N(_00047_),
    .Q(\dp.rf.rf[15][31] ));
 sg13g2_dfrbp_1 _16304_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_08518_),
    .D(_01278_),
    .Q_N(_00016_),
    .Q(\dp.rf.rf[16][0] ));
 sg13g2_dfrbp_1 _16305_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01279_),
    .Q_N(_01006_),
    .Q(\dp.rf.rf[16][1] ));
 sg13g2_dfrbp_1 _16306_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01280_),
    .Q_N(_00974_),
    .Q(\dp.rf.rf[16][2] ));
 sg13g2_dfrbp_1 _16307_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01281_),
    .Q_N(_00942_),
    .Q(\dp.rf.rf[16][3] ));
 sg13g2_dfrbp_1 _16308_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01282_),
    .Q_N(_00910_),
    .Q(\dp.rf.rf[16][4] ));
 sg13g2_dfrbp_1 _16309_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_08518_),
    .D(_01283_),
    .Q_N(_00878_),
    .Q(\dp.rf.rf[16][5] ));
 sg13g2_dfrbp_1 _16310_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01284_),
    .Q_N(_00846_),
    .Q(\dp.rf.rf[16][6] ));
 sg13g2_dfrbp_1 _16311_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01285_),
    .Q_N(_00814_),
    .Q(\dp.rf.rf[16][7] ));
 sg13g2_dfrbp_1 _16312_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01286_),
    .Q_N(_00782_),
    .Q(\dp.rf.rf[16][8] ));
 sg13g2_dfrbp_1 _16313_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01287_),
    .Q_N(_00750_),
    .Q(\dp.rf.rf[16][9] ));
 sg13g2_dfrbp_1 _16314_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_08518_),
    .D(_01288_),
    .Q_N(_00718_),
    .Q(\dp.rf.rf[16][10] ));
 sg13g2_dfrbp_1 _16315_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01289_),
    .Q_N(_00686_),
    .Q(\dp.rf.rf[16][11] ));
 sg13g2_dfrbp_1 _16316_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_08518_),
    .D(_01290_),
    .Q_N(_00654_),
    .Q(\dp.rf.rf[16][12] ));
 sg13g2_dfrbp_1 _16317_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_08518_),
    .D(_01291_),
    .Q_N(_00622_),
    .Q(\dp.rf.rf[16][13] ));
 sg13g2_dfrbp_1 _16318_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(_08518_),
    .D(_01292_),
    .Q_N(_00590_),
    .Q(\dp.rf.rf[16][14] ));
 sg13g2_dfrbp_1 _16319_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01293_),
    .Q_N(_00558_),
    .Q(\dp.rf.rf[16][15] ));
 sg13g2_dfrbp_1 _16320_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01294_),
    .Q_N(_00526_),
    .Q(\dp.rf.rf[16][16] ));
 sg13g2_dfrbp_1 _16321_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(_08518_),
    .D(_01295_),
    .Q_N(_00494_),
    .Q(\dp.rf.rf[16][17] ));
 sg13g2_dfrbp_1 _16322_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(_01296_),
    .Q_N(_00463_),
    .Q(\dp.rf.rf[16][18] ));
 sg13g2_dfrbp_1 _16323_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(_01297_),
    .Q_N(_00431_),
    .Q(\dp.rf.rf[16][19] ));
 sg13g2_dfrbp_1 _16324_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01298_),
    .Q_N(_00400_),
    .Q(\dp.rf.rf[16][20] ));
 sg13g2_dfrbp_1 _16325_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01299_),
    .Q_N(_00368_),
    .Q(\dp.rf.rf[16][21] ));
 sg13g2_dfrbp_1 _16326_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01300_),
    .Q_N(_00336_),
    .Q(\dp.rf.rf[16][22] ));
 sg13g2_dfrbp_1 _16327_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_08518_),
    .D(_01301_),
    .Q_N(_00304_),
    .Q(\dp.rf.rf[16][23] ));
 sg13g2_dfrbp_1 _16328_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(_08518_),
    .D(_01302_),
    .Q_N(_00272_),
    .Q(\dp.rf.rf[16][24] ));
 sg13g2_dfrbp_1 _16329_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01303_),
    .Q_N(_00240_),
    .Q(\dp.rf.rf[16][25] ));
 sg13g2_dfrbp_1 _16330_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01304_),
    .Q_N(_00208_),
    .Q(\dp.rf.rf[16][26] ));
 sg13g2_dfrbp_1 _16331_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01305_),
    .Q_N(_00176_),
    .Q(\dp.rf.rf[16][27] ));
 sg13g2_dfrbp_1 _16332_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01306_),
    .Q_N(_00144_),
    .Q(\dp.rf.rf[16][28] ));
 sg13g2_dfrbp_1 _16333_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01307_),
    .Q_N(_00112_),
    .Q(\dp.rf.rf[16][29] ));
 sg13g2_dfrbp_1 _16334_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01308_),
    .Q_N(_00080_),
    .Q(\dp.rf.rf[16][30] ));
 sg13g2_dfrbp_1 _16335_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01309_),
    .Q_N(_00048_),
    .Q(\dp.rf.rf[16][31] ));
 sg13g2_dfrbp_1 _16336_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_08518_),
    .D(_01310_),
    .Q_N(_00017_),
    .Q(\dp.rf.rf[17][0] ));
 sg13g2_dfrbp_1 _16337_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01311_),
    .Q_N(_01007_),
    .Q(\dp.rf.rf[17][1] ));
 sg13g2_dfrbp_1 _16338_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01312_),
    .Q_N(_00975_),
    .Q(\dp.rf.rf[17][2] ));
 sg13g2_dfrbp_1 _16339_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01313_),
    .Q_N(_00943_),
    .Q(\dp.rf.rf[17][3] ));
 sg13g2_dfrbp_1 _16340_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01314_),
    .Q_N(_00911_),
    .Q(\dp.rf.rf[17][4] ));
 sg13g2_dfrbp_1 _16341_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_08518_),
    .D(_01315_),
    .Q_N(_00879_),
    .Q(\dp.rf.rf[17][5] ));
 sg13g2_dfrbp_1 _16342_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01316_),
    .Q_N(_00847_),
    .Q(\dp.rf.rf[17][6] ));
 sg13g2_dfrbp_1 _16343_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01317_),
    .Q_N(_00815_),
    .Q(\dp.rf.rf[17][7] ));
 sg13g2_dfrbp_1 _16344_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01318_),
    .Q_N(_00783_),
    .Q(\dp.rf.rf[17][8] ));
 sg13g2_dfrbp_1 _16345_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01319_),
    .Q_N(_00751_),
    .Q(\dp.rf.rf[17][9] ));
 sg13g2_dfrbp_1 _16346_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01320_),
    .Q_N(_00719_),
    .Q(\dp.rf.rf[17][10] ));
 sg13g2_dfrbp_1 _16347_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01321_),
    .Q_N(_00687_),
    .Q(\dp.rf.rf[17][11] ));
 sg13g2_dfrbp_1 _16348_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_08518_),
    .D(_01322_),
    .Q_N(_00655_),
    .Q(\dp.rf.rf[17][12] ));
 sg13g2_dfrbp_1 _16349_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(_08518_),
    .D(_01323_),
    .Q_N(_00623_),
    .Q(\dp.rf.rf[17][13] ));
 sg13g2_dfrbp_1 _16350_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(_08518_),
    .D(_01324_),
    .Q_N(_00591_),
    .Q(\dp.rf.rf[17][14] ));
 sg13g2_dfrbp_1 _16351_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01325_),
    .Q_N(_00559_),
    .Q(\dp.rf.rf[17][15] ));
 sg13g2_dfrbp_1 _16352_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01326_),
    .Q_N(_00527_),
    .Q(\dp.rf.rf[17][16] ));
 sg13g2_dfrbp_1 _16353_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(_08518_),
    .D(_01327_),
    .Q_N(_00495_),
    .Q(\dp.rf.rf[17][17] ));
 sg13g2_dfrbp_1 _16354_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(_01328_),
    .Q_N(_00464_),
    .Q(\dp.rf.rf[17][18] ));
 sg13g2_dfrbp_1 _16355_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_01329_),
    .Q_N(_00432_),
    .Q(\dp.rf.rf[17][19] ));
 sg13g2_dfrbp_1 _16356_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01330_),
    .Q_N(_00401_),
    .Q(\dp.rf.rf[17][20] ));
 sg13g2_dfrbp_1 _16357_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01331_),
    .Q_N(_00369_),
    .Q(\dp.rf.rf[17][21] ));
 sg13g2_dfrbp_1 _16358_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(_08518_),
    .D(_01332_),
    .Q_N(_00337_),
    .Q(\dp.rf.rf[17][22] ));
 sg13g2_dfrbp_1 _16359_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_08518_),
    .D(_01333_),
    .Q_N(_00305_),
    .Q(\dp.rf.rf[17][23] ));
 sg13g2_dfrbp_1 _16360_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(_08518_),
    .D(_01334_),
    .Q_N(_00273_),
    .Q(\dp.rf.rf[17][24] ));
 sg13g2_dfrbp_1 _16361_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01335_),
    .Q_N(_00241_),
    .Q(\dp.rf.rf[17][25] ));
 sg13g2_dfrbp_1 _16362_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01336_),
    .Q_N(_00209_),
    .Q(\dp.rf.rf[17][26] ));
 sg13g2_dfrbp_1 _16363_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01337_),
    .Q_N(_00177_),
    .Q(\dp.rf.rf[17][27] ));
 sg13g2_dfrbp_1 _16364_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(_08518_),
    .D(_01338_),
    .Q_N(_00145_),
    .Q(\dp.rf.rf[17][28] ));
 sg13g2_dfrbp_1 _16365_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01339_),
    .Q_N(_00113_),
    .Q(\dp.rf.rf[17][29] ));
 sg13g2_dfrbp_1 _16366_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01340_),
    .Q_N(_00081_),
    .Q(\dp.rf.rf[17][30] ));
 sg13g2_dfrbp_1 _16367_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01341_),
    .Q_N(_00049_),
    .Q(\dp.rf.rf[17][31] ));
 sg13g2_dfrbp_1 _16368_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_08518_),
    .D(_01342_),
    .Q_N(_00018_),
    .Q(\dp.rf.rf[18][0] ));
 sg13g2_dfrbp_1 _16369_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01343_),
    .Q_N(_01008_),
    .Q(\dp.rf.rf[18][1] ));
 sg13g2_dfrbp_1 _16370_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01344_),
    .Q_N(_00976_),
    .Q(\dp.rf.rf[18][2] ));
 sg13g2_dfrbp_1 _16371_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01345_),
    .Q_N(_00944_),
    .Q(\dp.rf.rf[18][3] ));
 sg13g2_dfrbp_1 _16372_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01346_),
    .Q_N(_00912_),
    .Q(\dp.rf.rf[18][4] ));
 sg13g2_dfrbp_1 _16373_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_08518_),
    .D(_01347_),
    .Q_N(_00880_),
    .Q(\dp.rf.rf[18][5] ));
 sg13g2_dfrbp_1 _16374_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01348_),
    .Q_N(_00848_),
    .Q(\dp.rf.rf[18][6] ));
 sg13g2_dfrbp_1 _16375_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01349_),
    .Q_N(_00816_),
    .Q(\dp.rf.rf[18][7] ));
 sg13g2_dfrbp_1 _16376_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01350_),
    .Q_N(_00784_),
    .Q(\dp.rf.rf[18][8] ));
 sg13g2_dfrbp_1 _16377_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01351_),
    .Q_N(_00752_),
    .Q(\dp.rf.rf[18][9] ));
 sg13g2_dfrbp_1 _16378_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01352_),
    .Q_N(_00720_),
    .Q(\dp.rf.rf[18][10] ));
 sg13g2_dfrbp_1 _16379_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01353_),
    .Q_N(_00688_),
    .Q(\dp.rf.rf[18][11] ));
 sg13g2_dfrbp_1 _16380_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_08518_),
    .D(_01354_),
    .Q_N(_00656_),
    .Q(\dp.rf.rf[18][12] ));
 sg13g2_dfrbp_1 _16381_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_08518_),
    .D(_01355_),
    .Q_N(_00624_),
    .Q(\dp.rf.rf[18][13] ));
 sg13g2_dfrbp_1 _16382_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(_08518_),
    .D(_01356_),
    .Q_N(_00592_),
    .Q(\dp.rf.rf[18][14] ));
 sg13g2_dfrbp_1 _16383_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01357_),
    .Q_N(_00560_),
    .Q(\dp.rf.rf[18][15] ));
 sg13g2_dfrbp_1 _16384_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01358_),
    .Q_N(_00528_),
    .Q(\dp.rf.rf[18][16] ));
 sg13g2_dfrbp_1 _16385_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(_08518_),
    .D(_01359_),
    .Q_N(_00496_),
    .Q(\dp.rf.rf[18][17] ));
 sg13g2_dfrbp_1 _16386_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01360_),
    .Q_N(_00465_),
    .Q(\dp.rf.rf[18][18] ));
 sg13g2_dfrbp_1 _16387_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(_01361_),
    .Q_N(_00433_),
    .Q(\dp.rf.rf[18][19] ));
 sg13g2_dfrbp_1 _16388_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01362_),
    .Q_N(_00402_),
    .Q(\dp.rf.rf[18][20] ));
 sg13g2_dfrbp_1 _16389_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01363_),
    .Q_N(_00370_),
    .Q(\dp.rf.rf[18][21] ));
 sg13g2_dfrbp_1 _16390_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(_08518_),
    .D(_01364_),
    .Q_N(_00338_),
    .Q(\dp.rf.rf[18][22] ));
 sg13g2_dfrbp_1 _16391_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_01365_),
    .Q_N(_00306_),
    .Q(\dp.rf.rf[18][23] ));
 sg13g2_dfrbp_1 _16392_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(_08518_),
    .D(_01366_),
    .Q_N(_00274_),
    .Q(\dp.rf.rf[18][24] ));
 sg13g2_dfrbp_1 _16393_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01367_),
    .Q_N(_00242_),
    .Q(\dp.rf.rf[18][25] ));
 sg13g2_dfrbp_1 _16394_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01368_),
    .Q_N(_00210_),
    .Q(\dp.rf.rf[18][26] ));
 sg13g2_dfrbp_1 _16395_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01369_),
    .Q_N(_00178_),
    .Q(\dp.rf.rf[18][27] ));
 sg13g2_dfrbp_1 _16396_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01370_),
    .Q_N(_00146_),
    .Q(\dp.rf.rf[18][28] ));
 sg13g2_dfrbp_1 _16397_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01371_),
    .Q_N(_00114_),
    .Q(\dp.rf.rf[18][29] ));
 sg13g2_dfrbp_1 _16398_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01372_),
    .Q_N(_00082_),
    .Q(\dp.rf.rf[18][30] ));
 sg13g2_dfrbp_1 _16399_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01373_),
    .Q_N(_00050_),
    .Q(\dp.rf.rf[18][31] ));
 sg13g2_dfrbp_1 _16400_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_08518_),
    .D(_01374_),
    .Q_N(_00001_),
    .Q(\dp.rf.rf[1][0] ));
 sg13g2_dfrbp_1 _16401_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_08518_),
    .D(_01375_),
    .Q_N(_00991_),
    .Q(\dp.rf.rf[1][1] ));
 sg13g2_dfrbp_1 _16402_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01376_),
    .Q_N(_00959_),
    .Q(\dp.rf.rf[1][2] ));
 sg13g2_dfrbp_1 _16403_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01377_),
    .Q_N(_00927_),
    .Q(\dp.rf.rf[1][3] ));
 sg13g2_dfrbp_1 _16404_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_01378_),
    .Q_N(_00895_),
    .Q(\dp.rf.rf[1][4] ));
 sg13g2_dfrbp_1 _16405_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_08518_),
    .D(_01379_),
    .Q_N(_00863_),
    .Q(\dp.rf.rf[1][5] ));
 sg13g2_dfrbp_1 _16406_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_08518_),
    .D(_01380_),
    .Q_N(_00831_),
    .Q(\dp.rf.rf[1][6] ));
 sg13g2_dfrbp_1 _16407_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01381_),
    .Q_N(_00799_),
    .Q(\dp.rf.rf[1][7] ));
 sg13g2_dfrbp_1 _16408_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_01382_),
    .Q_N(_00767_),
    .Q(\dp.rf.rf[1][8] ));
 sg13g2_dfrbp_1 _16409_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_01383_),
    .Q_N(_00735_),
    .Q(\dp.rf.rf[1][9] ));
 sg13g2_dfrbp_1 _16410_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01384_),
    .Q_N(_00703_),
    .Q(\dp.rf.rf[1][10] ));
 sg13g2_dfrbp_1 _16411_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01385_),
    .Q_N(_00671_),
    .Q(\dp.rf.rf[1][11] ));
 sg13g2_dfrbp_1 _16412_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_08518_),
    .D(_01386_),
    .Q_N(_00639_),
    .Q(\dp.rf.rf[1][12] ));
 sg13g2_dfrbp_1 _16413_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01387_),
    .Q_N(_00607_),
    .Q(\dp.rf.rf[1][13] ));
 sg13g2_dfrbp_1 _16414_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(_01388_),
    .Q_N(_00575_),
    .Q(\dp.rf.rf[1][14] ));
 sg13g2_dfrbp_1 _16415_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_08518_),
    .D(_01389_),
    .Q_N(_00543_),
    .Q(\dp.rf.rf[1][15] ));
 sg13g2_dfrbp_1 _16416_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_08518_),
    .D(_01390_),
    .Q_N(_00511_),
    .Q(\dp.rf.rf[1][16] ));
 sg13g2_dfrbp_1 _16417_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(_08518_),
    .D(_01391_),
    .Q_N(_00479_),
    .Q(\dp.rf.rf[1][17] ));
 sg13g2_dfrbp_1 _16418_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01392_),
    .Q_N(_00448_),
    .Q(\dp.rf.rf[1][18] ));
 sg13g2_dfrbp_1 _16419_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_01393_),
    .Q_N(_00416_),
    .Q(\dp.rf.rf[1][19] ));
 sg13g2_dfrbp_1 _16420_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(_08518_),
    .D(_01394_),
    .Q_N(_00385_),
    .Q(\dp.rf.rf[1][20] ));
 sg13g2_dfrbp_1 _16421_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01395_),
    .Q_N(_00353_),
    .Q(\dp.rf.rf[1][21] ));
 sg13g2_dfrbp_1 _16422_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(_08518_),
    .D(_01396_),
    .Q_N(_00321_),
    .Q(\dp.rf.rf[1][22] ));
 sg13g2_dfrbp_1 _16423_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01397_),
    .Q_N(_00289_),
    .Q(\dp.rf.rf[1][23] ));
 sg13g2_dfrbp_1 _16424_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(_08518_),
    .D(_01398_),
    .Q_N(_00257_),
    .Q(\dp.rf.rf[1][24] ));
 sg13g2_dfrbp_1 _16425_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01399_),
    .Q_N(_00225_),
    .Q(\dp.rf.rf[1][25] ));
 sg13g2_dfrbp_1 _16426_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(_08518_),
    .D(_01400_),
    .Q_N(_00193_),
    .Q(\dp.rf.rf[1][26] ));
 sg13g2_dfrbp_1 _16427_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01401_),
    .Q_N(_00161_),
    .Q(\dp.rf.rf[1][27] ));
 sg13g2_dfrbp_1 _16428_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01402_),
    .Q_N(_00129_),
    .Q(\dp.rf.rf[1][28] ));
 sg13g2_dfrbp_1 _16429_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01403_),
    .Q_N(_00097_),
    .Q(\dp.rf.rf[1][29] ));
 sg13g2_dfrbp_1 _16430_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01404_),
    .Q_N(_00065_),
    .Q(\dp.rf.rf[1][30] ));
 sg13g2_dfrbp_1 _16431_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_08518_),
    .D(_01405_),
    .Q_N(_00033_),
    .Q(\dp.rf.rf[1][31] ));
 sg13g2_dfrbp_1 _16432_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_08518_),
    .D(_01406_),
    .Q_N(_00020_),
    .Q(\dp.rf.rf[20][0] ));
 sg13g2_dfrbp_1 _16433_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01407_),
    .Q_N(_01010_),
    .Q(\dp.rf.rf[20][1] ));
 sg13g2_dfrbp_1 _16434_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01408_),
    .Q_N(_00978_),
    .Q(\dp.rf.rf[20][2] ));
 sg13g2_dfrbp_1 _16435_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_01409_),
    .Q_N(_00946_),
    .Q(\dp.rf.rf[20][3] ));
 sg13g2_dfrbp_1 _16436_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(_01410_),
    .Q_N(_00914_),
    .Q(\dp.rf.rf[20][4] ));
 sg13g2_dfrbp_1 _16437_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_08518_),
    .D(_01411_),
    .Q_N(_00882_),
    .Q(\dp.rf.rf[20][5] ));
 sg13g2_dfrbp_1 _16438_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01412_),
    .Q_N(_00850_),
    .Q(\dp.rf.rf[20][6] ));
 sg13g2_dfrbp_1 _16439_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01413_),
    .Q_N(_00818_),
    .Q(\dp.rf.rf[20][7] ));
 sg13g2_dfrbp_1 _16440_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_01414_),
    .Q_N(_00786_),
    .Q(\dp.rf.rf[20][8] ));
 sg13g2_dfrbp_1 _16441_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(_01415_),
    .Q_N(_00754_),
    .Q(\dp.rf.rf[20][9] ));
 sg13g2_dfrbp_1 _16442_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01416_),
    .Q_N(_00722_),
    .Q(\dp.rf.rf[20][10] ));
 sg13g2_dfrbp_1 _16443_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_01417_),
    .Q_N(_00690_),
    .Q(\dp.rf.rf[20][11] ));
 sg13g2_dfrbp_1 _16444_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01418_),
    .Q_N(_00658_),
    .Q(\dp.rf.rf[20][12] ));
 sg13g2_dfrbp_1 _16445_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_08518_),
    .D(_01419_),
    .Q_N(_00626_),
    .Q(\dp.rf.rf[20][13] ));
 sg13g2_dfrbp_1 _16446_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01420_),
    .Q_N(_00594_),
    .Q(\dp.rf.rf[20][14] ));
 sg13g2_dfrbp_1 _16447_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01421_),
    .Q_N(_00562_),
    .Q(\dp.rf.rf[20][15] ));
 sg13g2_dfrbp_1 _16448_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_08518_),
    .D(_01422_),
    .Q_N(_00530_),
    .Q(\dp.rf.rf[20][16] ));
 sg13g2_dfrbp_1 _16449_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01423_),
    .Q_N(_00498_),
    .Q(\dp.rf.rf[20][17] ));
 sg13g2_dfrbp_1 _16450_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_01424_),
    .Q_N(_00467_),
    .Q(\dp.rf.rf[20][18] ));
 sg13g2_dfrbp_1 _16451_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01425_),
    .Q_N(_00435_),
    .Q(\dp.rf.rf[20][19] ));
 sg13g2_dfrbp_1 _16452_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01426_),
    .Q_N(_00404_),
    .Q(\dp.rf.rf[20][20] ));
 sg13g2_dfrbp_1 _16453_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01427_),
    .Q_N(_00372_),
    .Q(\dp.rf.rf[20][21] ));
 sg13g2_dfrbp_1 _16454_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01428_),
    .Q_N(_00340_),
    .Q(\dp.rf.rf[20][22] ));
 sg13g2_dfrbp_1 _16455_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01429_),
    .Q_N(_00308_),
    .Q(\dp.rf.rf[20][23] ));
 sg13g2_dfrbp_1 _16456_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01430_),
    .Q_N(_00276_),
    .Q(\dp.rf.rf[20][24] ));
 sg13g2_dfrbp_1 _16457_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01431_),
    .Q_N(_00244_),
    .Q(\dp.rf.rf[20][25] ));
 sg13g2_dfrbp_1 _16458_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01432_),
    .Q_N(_00212_),
    .Q(\dp.rf.rf[20][26] ));
 sg13g2_dfrbp_1 _16459_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(_08518_),
    .D(_01433_),
    .Q_N(_00180_),
    .Q(\dp.rf.rf[20][27] ));
 sg13g2_dfrbp_1 _16460_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01434_),
    .Q_N(_00148_),
    .Q(\dp.rf.rf[20][28] ));
 sg13g2_dfrbp_1 _16461_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01435_),
    .Q_N(_00116_),
    .Q(\dp.rf.rf[20][29] ));
 sg13g2_dfrbp_1 _16462_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01436_),
    .Q_N(_00084_),
    .Q(\dp.rf.rf[20][30] ));
 sg13g2_dfrbp_1 _16463_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01437_),
    .Q_N(_00052_),
    .Q(\dp.rf.rf[20][31] ));
 sg13g2_dfrbp_1 _16464_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01438_),
    .Q_N(_00008_),
    .Q(\dp.rf.rf[8][0] ));
 sg13g2_dfrbp_1 _16465_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01439_),
    .Q_N(_00998_),
    .Q(\dp.rf.rf[8][1] ));
 sg13g2_dfrbp_1 _16466_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01440_),
    .Q_N(_00966_),
    .Q(\dp.rf.rf[8][2] ));
 sg13g2_dfrbp_1 _16467_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(_08518_),
    .D(_01441_),
    .Q_N(_00934_),
    .Q(\dp.rf.rf[8][3] ));
 sg13g2_dfrbp_1 _16468_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_08518_),
    .D(_01442_),
    .Q_N(_00902_),
    .Q(\dp.rf.rf[8][4] ));
 sg13g2_dfrbp_1 _16469_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_08518_),
    .D(_01443_),
    .Q_N(_00870_),
    .Q(\dp.rf.rf[8][5] ));
 sg13g2_dfrbp_1 _16470_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_08518_),
    .D(_01444_),
    .Q_N(_00838_),
    .Q(\dp.rf.rf[8][6] ));
 sg13g2_dfrbp_1 _16471_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_01445_),
    .Q_N(_00806_),
    .Q(\dp.rf.rf[8][7] ));
 sg13g2_dfrbp_1 _16472_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_08518_),
    .D(_01446_),
    .Q_N(_00774_),
    .Q(\dp.rf.rf[8][8] ));
 sg13g2_dfrbp_1 _16473_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01447_),
    .Q_N(_00742_),
    .Q(\dp.rf.rf[8][9] ));
 sg13g2_dfrbp_1 _16474_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01448_),
    .Q_N(_00710_),
    .Q(\dp.rf.rf[8][10] ));
 sg13g2_dfrbp_1 _16475_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01449_),
    .Q_N(_00678_),
    .Q(\dp.rf.rf[8][11] ));
 sg13g2_dfrbp_1 _16476_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01450_),
    .Q_N(_00646_),
    .Q(\dp.rf.rf[8][12] ));
 sg13g2_dfrbp_1 _16477_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_08518_),
    .D(_01451_),
    .Q_N(_00614_),
    .Q(\dp.rf.rf[8][13] ));
 sg13g2_dfrbp_1 _16478_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01452_),
    .Q_N(_00582_),
    .Q(\dp.rf.rf[8][14] ));
 sg13g2_dfrbp_1 _16479_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_08518_),
    .D(_01453_),
    .Q_N(_00550_),
    .Q(\dp.rf.rf[8][15] ));
 sg13g2_dfrbp_1 _16480_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_01454_),
    .Q_N(_00518_),
    .Q(\dp.rf.rf[8][16] ));
 sg13g2_dfrbp_1 _16481_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(_08518_),
    .D(_01455_),
    .Q_N(_00486_),
    .Q(\dp.rf.rf[8][17] ));
 sg13g2_dfrbp_1 _16482_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(_01456_),
    .Q_N(_00455_),
    .Q(\dp.rf.rf[8][18] ));
 sg13g2_dfrbp_1 _16483_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(_01457_),
    .Q_N(_00423_),
    .Q(\dp.rf.rf[8][19] ));
 sg13g2_dfrbp_1 _16484_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(_08518_),
    .D(_01458_),
    .Q_N(_00392_),
    .Q(\dp.rf.rf[8][20] ));
 sg13g2_dfrbp_1 _16485_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01459_),
    .Q_N(_00360_),
    .Q(\dp.rf.rf[8][21] ));
 sg13g2_dfrbp_1 _16486_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01460_),
    .Q_N(_00328_),
    .Q(\dp.rf.rf[8][22] ));
 sg13g2_dfrbp_1 _16487_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01461_),
    .Q_N(_00296_),
    .Q(\dp.rf.rf[8][23] ));
 sg13g2_dfrbp_1 _16488_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(_08518_),
    .D(_01462_),
    .Q_N(_00264_),
    .Q(\dp.rf.rf[8][24] ));
 sg13g2_dfrbp_1 _16489_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01463_),
    .Q_N(_00232_),
    .Q(\dp.rf.rf[8][25] ));
 sg13g2_dfrbp_1 _16490_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01464_),
    .Q_N(_00200_),
    .Q(\dp.rf.rf[8][26] ));
 sg13g2_dfrbp_1 _16491_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_01465_),
    .Q_N(_00168_),
    .Q(\dp.rf.rf[8][27] ));
 sg13g2_dfrbp_1 _16492_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01466_),
    .Q_N(_00136_),
    .Q(\dp.rf.rf[8][28] ));
 sg13g2_dfrbp_1 _16493_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01467_),
    .Q_N(_00104_),
    .Q(\dp.rf.rf[8][29] ));
 sg13g2_dfrbp_1 _16494_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01468_),
    .Q_N(_00072_),
    .Q(\dp.rf.rf[8][30] ));
 sg13g2_dfrbp_1 _16495_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_08518_),
    .D(_01469_),
    .Q_N(_00040_),
    .Q(\dp.rf.rf[8][31] ));
 sg13g2_dfrbp_1 _16496_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_08518_),
    .D(_01470_),
    .Q_N(_00010_),
    .Q(\dp.rf.rf[10][0] ));
 sg13g2_dfrbp_1 _16497_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01471_),
    .Q_N(_01000_),
    .Q(\dp.rf.rf[10][1] ));
 sg13g2_dfrbp_1 _16498_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01472_),
    .Q_N(_00968_),
    .Q(\dp.rf.rf[10][2] ));
 sg13g2_dfrbp_1 _16499_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(_08518_),
    .D(_01473_),
    .Q_N(_00936_),
    .Q(\dp.rf.rf[10][3] ));
 sg13g2_dfrbp_1 _16500_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_08518_),
    .D(_01474_),
    .Q_N(_00904_),
    .Q(\dp.rf.rf[10][4] ));
 sg13g2_dfrbp_1 _16501_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_08518_),
    .D(_01475_),
    .Q_N(_00872_),
    .Q(\dp.rf.rf[10][5] ));
 sg13g2_dfrbp_1 _16502_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_08518_),
    .D(_01476_),
    .Q_N(_00840_),
    .Q(\dp.rf.rf[10][6] ));
 sg13g2_dfrbp_1 _16503_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_01477_),
    .Q_N(_00808_),
    .Q(\dp.rf.rf[10][7] ));
 sg13g2_dfrbp_1 _16504_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_01478_),
    .Q_N(_00776_),
    .Q(\dp.rf.rf[10][8] ));
 sg13g2_dfrbp_1 _16505_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01479_),
    .Q_N(_00744_),
    .Q(\dp.rf.rf[10][9] ));
 sg13g2_dfrbp_1 _16506_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01480_),
    .Q_N(_00712_),
    .Q(\dp.rf.rf[10][10] ));
 sg13g2_dfrbp_1 _16507_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01481_),
    .Q_N(_00680_),
    .Q(\dp.rf.rf[10][11] ));
 sg13g2_dfrbp_1 _16508_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01482_),
    .Q_N(_00648_),
    .Q(\dp.rf.rf[10][12] ));
 sg13g2_dfrbp_1 _16509_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_08518_),
    .D(_01483_),
    .Q_N(_00616_),
    .Q(\dp.rf.rf[10][13] ));
 sg13g2_dfrbp_1 _16510_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01484_),
    .Q_N(_00584_),
    .Q(\dp.rf.rf[10][14] ));
 sg13g2_dfrbp_1 _16511_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_01485_),
    .Q_N(_00552_),
    .Q(\dp.rf.rf[10][15] ));
 sg13g2_dfrbp_1 _16512_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_01486_),
    .Q_N(_00520_),
    .Q(\dp.rf.rf[10][16] ));
 sg13g2_dfrbp_1 _16513_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(_08518_),
    .D(_01487_),
    .Q_N(_00488_),
    .Q(\dp.rf.rf[10][17] ));
 sg13g2_dfrbp_1 _16514_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(_01488_),
    .Q_N(_00457_),
    .Q(\dp.rf.rf[10][18] ));
 sg13g2_dfrbp_1 _16515_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(_01489_),
    .Q_N(_00425_),
    .Q(\dp.rf.rf[10][19] ));
 sg13g2_dfrbp_1 _16516_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(_08518_),
    .D(_01490_),
    .Q_N(_00394_),
    .Q(\dp.rf.rf[10][20] ));
 sg13g2_dfrbp_1 _16517_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01491_),
    .Q_N(_00362_),
    .Q(\dp.rf.rf[10][21] ));
 sg13g2_dfrbp_1 _16518_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01492_),
    .Q_N(_00330_),
    .Q(\dp.rf.rf[10][22] ));
 sg13g2_dfrbp_1 _16519_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01493_),
    .Q_N(_00298_),
    .Q(\dp.rf.rf[10][23] ));
 sg13g2_dfrbp_1 _16520_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01494_),
    .Q_N(_00266_),
    .Q(\dp.rf.rf[10][24] ));
 sg13g2_dfrbp_1 _16521_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01495_),
    .Q_N(_00234_),
    .Q(\dp.rf.rf[10][25] ));
 sg13g2_dfrbp_1 _16522_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01496_),
    .Q_N(_00202_),
    .Q(\dp.rf.rf[10][26] ));
 sg13g2_dfrbp_1 _16523_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_01497_),
    .Q_N(_00170_),
    .Q(\dp.rf.rf[10][27] ));
 sg13g2_dfrbp_1 _16524_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01498_),
    .Q_N(_00138_),
    .Q(\dp.rf.rf[10][28] ));
 sg13g2_dfrbp_1 _16525_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01499_),
    .Q_N(_00106_),
    .Q(\dp.rf.rf[10][29] ));
 sg13g2_dfrbp_1 _16526_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01500_),
    .Q_N(_00074_),
    .Q(\dp.rf.rf[10][30] ));
 sg13g2_dfrbp_1 _16527_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_01501_),
    .Q_N(_00042_),
    .Q(\dp.rf.rf[10][31] ));
 sg13g2_dfrbp_1 _16528_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_08518_),
    .D(_01502_),
    .Q_N(_00007_),
    .Q(\dp.rf.rf[7][0] ));
 sg13g2_dfrbp_1 _16529_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01503_),
    .Q_N(_00997_),
    .Q(\dp.rf.rf[7][1] ));
 sg13g2_dfrbp_1 _16530_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01504_),
    .Q_N(_00965_),
    .Q(\dp.rf.rf[7][2] ));
 sg13g2_dfrbp_1 _16531_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(_08518_),
    .D(_01505_),
    .Q_N(_00933_),
    .Q(\dp.rf.rf[7][3] ));
 sg13g2_dfrbp_1 _16532_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(_01506_),
    .Q_N(_00901_),
    .Q(\dp.rf.rf[7][4] ));
 sg13g2_dfrbp_1 _16533_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_08518_),
    .D(_01507_),
    .Q_N(_00869_),
    .Q(\dp.rf.rf[7][5] ));
 sg13g2_dfrbp_1 _16534_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_01508_),
    .Q_N(_00837_),
    .Q(\dp.rf.rf[7][6] ));
 sg13g2_dfrbp_1 _16535_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01509_),
    .Q_N(_00805_),
    .Q(\dp.rf.rf[7][7] ));
 sg13g2_dfrbp_1 _16536_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01510_),
    .Q_N(_00773_),
    .Q(\dp.rf.rf[7][8] ));
 sg13g2_dfrbp_1 _16537_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_01511_),
    .Q_N(_00741_),
    .Q(\dp.rf.rf[7][9] ));
 sg13g2_dfrbp_1 _16538_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01512_),
    .Q_N(_00709_),
    .Q(\dp.rf.rf[7][10] ));
 sg13g2_dfrbp_1 _16539_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_01513_),
    .Q_N(_00677_),
    .Q(\dp.rf.rf[7][11] ));
 sg13g2_dfrbp_1 _16540_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01514_),
    .Q_N(_00645_),
    .Q(\dp.rf.rf[7][12] ));
 sg13g2_dfrbp_1 _16541_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_08518_),
    .D(_01515_),
    .Q_N(_00613_),
    .Q(\dp.rf.rf[7][13] ));
 sg13g2_dfrbp_1 _16542_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(_08518_),
    .D(_01516_),
    .Q_N(_00581_),
    .Q(\dp.rf.rf[7][14] ));
 sg13g2_dfrbp_1 _16543_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_01517_),
    .Q_N(_00549_),
    .Q(\dp.rf.rf[7][15] ));
 sg13g2_dfrbp_1 _16544_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_08518_),
    .D(_01518_),
    .Q_N(_00517_),
    .Q(\dp.rf.rf[7][16] ));
 sg13g2_dfrbp_1 _16545_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(_08518_),
    .D(_01519_),
    .Q_N(_00485_),
    .Q(\dp.rf.rf[7][17] ));
 sg13g2_dfrbp_1 _16546_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(_01520_),
    .Q_N(_00454_),
    .Q(\dp.rf.rf[7][18] ));
 sg13g2_dfrbp_1 _16547_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_01521_),
    .Q_N(_00422_),
    .Q(\dp.rf.rf[7][19] ));
 sg13g2_dfrbp_1 _16548_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01522_),
    .Q_N(_00391_),
    .Q(\dp.rf.rf[7][20] ));
 sg13g2_dfrbp_1 _16549_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01523_),
    .Q_N(_00359_),
    .Q(\dp.rf.rf[7][21] ));
 sg13g2_dfrbp_1 _16550_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(_08518_),
    .D(_01524_),
    .Q_N(_00327_),
    .Q(\dp.rf.rf[7][22] ));
 sg13g2_dfrbp_1 _16551_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_08518_),
    .D(_01525_),
    .Q_N(_00295_),
    .Q(\dp.rf.rf[7][23] ));
 sg13g2_dfrbp_1 _16552_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01526_),
    .Q_N(_00263_),
    .Q(\dp.rf.rf[7][24] ));
 sg13g2_dfrbp_1 _16553_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01527_),
    .Q_N(_00231_),
    .Q(\dp.rf.rf[7][25] ));
 sg13g2_dfrbp_1 _16554_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01528_),
    .Q_N(_00199_),
    .Q(\dp.rf.rf[7][26] ));
 sg13g2_dfrbp_1 _16555_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01529_),
    .Q_N(_00167_),
    .Q(\dp.rf.rf[7][27] ));
 sg13g2_dfrbp_1 _16556_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_01530_),
    .Q_N(_00135_),
    .Q(\dp.rf.rf[7][28] ));
 sg13g2_dfrbp_1 _16557_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01531_),
    .Q_N(_00103_),
    .Q(\dp.rf.rf[7][29] ));
 sg13g2_dfrbp_1 _16558_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01532_),
    .Q_N(_00071_),
    .Q(\dp.rf.rf[7][30] ));
 sg13g2_dfrbp_1 _16559_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01533_),
    .Q_N(_00039_),
    .Q(\dp.rf.rf[7][31] ));
 sg13g2_dfrbp_1 _16560_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][0] ),
    .Q_N(_00000_),
    .Q(\dp.rf.rf[0][0] ));
 sg13g2_dfrbp_1 _16561_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][1] ),
    .Q_N(_00990_),
    .Q(\dp.rf.rf[0][1] ));
 sg13g2_dfrbp_1 _16562_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][2] ),
    .Q_N(_00958_),
    .Q(\dp.rf.rf[0][2] ));
 sg13g2_dfrbp_1 _16563_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][3] ),
    .Q_N(_00926_),
    .Q(\dp.rf.rf[0][3] ));
 sg13g2_dfrbp_1 _16564_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][4] ),
    .Q_N(_00894_),
    .Q(\dp.rf.rf[0][4] ));
 sg13g2_dfrbp_1 _16565_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][5] ),
    .Q_N(_00862_),
    .Q(\dp.rf.rf[0][5] ));
 sg13g2_dfrbp_1 _16566_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][6] ),
    .Q_N(_00830_),
    .Q(\dp.rf.rf[0][6] ));
 sg13g2_dfrbp_1 _16567_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][7] ),
    .Q_N(_00798_),
    .Q(\dp.rf.rf[0][7] ));
 sg13g2_dfrbp_1 _16568_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][8] ),
    .Q_N(_00766_),
    .Q(\dp.rf.rf[0][8] ));
 sg13g2_dfrbp_1 _16569_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][9] ),
    .Q_N(_00734_),
    .Q(\dp.rf.rf[0][9] ));
 sg13g2_dfrbp_1 _16570_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][10] ),
    .Q_N(_00702_),
    .Q(\dp.rf.rf[0][10] ));
 sg13g2_dfrbp_1 _16571_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][11] ),
    .Q_N(_00670_),
    .Q(\dp.rf.rf[0][11] ));
 sg13g2_dfrbp_1 _16572_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][12] ),
    .Q_N(_00638_),
    .Q(\dp.rf.rf[0][12] ));
 sg13g2_dfrbp_1 _16573_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][13] ),
    .Q_N(_00606_),
    .Q(\dp.rf.rf[0][13] ));
 sg13g2_dfrbp_1 _16574_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][14] ),
    .Q_N(_00574_),
    .Q(\dp.rf.rf[0][14] ));
 sg13g2_dfrbp_1 _16575_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][15] ),
    .Q_N(_00542_),
    .Q(\dp.rf.rf[0][15] ));
 sg13g2_dfrbp_1 _16576_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][16] ),
    .Q_N(_00510_),
    .Q(\dp.rf.rf[0][16] ));
 sg13g2_dfrbp_1 _16577_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][18] ),
    .Q_N(_00447_),
    .Q(\dp.rf.rf[0][18] ));
 sg13g2_dfrbp_1 _16578_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][20] ),
    .Q_N(_00384_),
    .Q(\dp.rf.rf[0][20] ));
 sg13g2_dfrbp_1 _16579_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][21] ),
    .Q_N(_00352_),
    .Q(\dp.rf.rf[0][21] ));
 sg13g2_dfrbp_1 _16580_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][22] ),
    .Q_N(_00320_),
    .Q(\dp.rf.rf[0][22] ));
 sg13g2_dfrbp_1 _16581_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][23] ),
    .Q_N(_00288_),
    .Q(\dp.rf.rf[0][23] ));
 sg13g2_dfrbp_1 _16582_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][24] ),
    .Q_N(_00256_),
    .Q(\dp.rf.rf[0][24] ));
 sg13g2_dfrbp_1 _16583_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][25] ),
    .Q_N(_00224_),
    .Q(\dp.rf.rf[0][25] ));
 sg13g2_dfrbp_1 _16584_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][26] ),
    .Q_N(_00192_),
    .Q(\dp.rf.rf[0][26] ));
 sg13g2_dfrbp_1 _16585_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][27] ),
    .Q_N(_00160_),
    .Q(\dp.rf.rf[0][27] ));
 sg13g2_dfrbp_1 _16586_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][28] ),
    .Q_N(_00128_),
    .Q(\dp.rf.rf[0][28] ));
 sg13g2_dfrbp_1 _16587_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][29] ),
    .Q_N(_00096_),
    .Q(\dp.rf.rf[0][29] ));
 sg13g2_dfrbp_1 _16588_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][30] ),
    .Q_N(_00064_),
    .Q(\dp.rf.rf[0][30] ));
 sg13g2_dfrbp_1 _16589_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(\dp.rf.rf[0][31] ),
    .Q_N(_00032_),
    .Q(\dp.rf.rf[0][31] ));
 sg13g2_dfrbp_1 _16590_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_08518_),
    .D(_01564_),
    .Q_N(_00004_),
    .Q(\dp.rf.rf[4][0] ));
 sg13g2_dfrbp_1 _16591_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_08518_),
    .D(_01565_),
    .Q_N(_00994_),
    .Q(\dp.rf.rf[4][1] ));
 sg13g2_dfrbp_1 _16592_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01566_),
    .Q_N(_00962_),
    .Q(\dp.rf.rf[4][2] ));
 sg13g2_dfrbp_1 _16593_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(_08518_),
    .D(_01567_),
    .Q_N(_00930_),
    .Q(\dp.rf.rf[4][3] ));
 sg13g2_dfrbp_1 _16594_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(_01568_),
    .Q_N(_00898_),
    .Q(\dp.rf.rf[4][4] ));
 sg13g2_dfrbp_1 _16595_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_08518_),
    .D(_01569_),
    .Q_N(_00866_),
    .Q(\dp.rf.rf[4][5] ));
 sg13g2_dfrbp_1 _16596_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_08518_),
    .D(_01570_),
    .Q_N(_00834_),
    .Q(\dp.rf.rf[4][6] ));
 sg13g2_dfrbp_1 _16597_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01571_),
    .Q_N(_00802_),
    .Q(\dp.rf.rf[4][7] ));
 sg13g2_dfrbp_1 _16598_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01572_),
    .Q_N(_00770_),
    .Q(\dp.rf.rf[4][8] ));
 sg13g2_dfrbp_1 _16599_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_01573_),
    .Q_N(_00738_),
    .Q(\dp.rf.rf[4][9] ));
 sg13g2_dfrbp_1 _16600_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_08518_),
    .D(_01574_),
    .Q_N(_00706_),
    .Q(\dp.rf.rf[4][10] ));
 sg13g2_dfrbp_1 _16601_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_01575_),
    .Q_N(_00674_),
    .Q(\dp.rf.rf[4][11] ));
 sg13g2_dfrbp_1 _16602_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_08518_),
    .D(_01576_),
    .Q_N(_00642_),
    .Q(\dp.rf.rf[4][12] ));
 sg13g2_dfrbp_1 _16603_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_01577_),
    .Q_N(_00610_),
    .Q(\dp.rf.rf[4][13] ));
 sg13g2_dfrbp_1 _16604_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01578_),
    .Q_N(_00578_),
    .Q(\dp.rf.rf[4][14] ));
 sg13g2_dfrbp_1 _16605_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_01579_),
    .Q_N(_00546_),
    .Q(\dp.rf.rf[4][15] ));
 sg13g2_dfrbp_1 _16606_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_01580_),
    .Q_N(_00514_),
    .Q(\dp.rf.rf[4][16] ));
 sg13g2_dfrbp_1 _16607_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(_08518_),
    .D(_01581_),
    .Q_N(_00482_),
    .Q(\dp.rf.rf[4][17] ));
 sg13g2_dfrbp_1 _16608_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_01582_),
    .Q_N(_00451_),
    .Q(\dp.rf.rf[4][18] ));
 sg13g2_dfrbp_1 _16609_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_01583_),
    .Q_N(_00419_),
    .Q(\dp.rf.rf[4][19] ));
 sg13g2_dfrbp_1 _16610_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01584_),
    .Q_N(_00388_),
    .Q(\dp.rf.rf[4][20] ));
 sg13g2_dfrbp_1 _16611_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01585_),
    .Q_N(_00356_),
    .Q(\dp.rf.rf[4][21] ));
 sg13g2_dfrbp_1 _16612_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(_08518_),
    .D(_01586_),
    .Q_N(_00324_),
    .Q(\dp.rf.rf[4][22] ));
 sg13g2_dfrbp_1 _16613_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_01587_),
    .Q_N(_00292_),
    .Q(\dp.rf.rf[4][23] ));
 sg13g2_dfrbp_1 _16614_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01588_),
    .Q_N(_00260_),
    .Q(\dp.rf.rf[4][24] ));
 sg13g2_dfrbp_1 _16615_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01589_),
    .Q_N(_00228_),
    .Q(\dp.rf.rf[4][25] ));
 sg13g2_dfrbp_1 _16616_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01590_),
    .Q_N(_00196_),
    .Q(\dp.rf.rf[4][26] ));
 sg13g2_dfrbp_1 _16617_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01591_),
    .Q_N(_00164_),
    .Q(\dp.rf.rf[4][27] ));
 sg13g2_dfrbp_1 _16618_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_01592_),
    .Q_N(_00132_),
    .Q(\dp.rf.rf[4][28] ));
 sg13g2_dfrbp_1 _16619_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01593_),
    .Q_N(_00100_),
    .Q(\dp.rf.rf[4][29] ));
 sg13g2_dfrbp_1 _16620_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01594_),
    .Q_N(_00068_),
    .Q(\dp.rf.rf[4][30] ));
 sg13g2_dfrbp_1 _16621_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01595_),
    .Q_N(_00036_),
    .Q(\dp.rf.rf[4][31] ));
 sg13g2_dfrbp_1 _16622_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net955),
    .D(\dp.ISRmux.d0[2] ),
    .Q_N(_01024_),
    .Q(net122));
 sg13g2_dfrbp_1 _16623_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net955),
    .D(\dp.ISRmux.d0[3] ),
    .Q_N(_01025_),
    .Q(net125));
 sg13g2_dfrbp_1 _16624_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net955),
    .D(\dp.ISRmux.d0[4] ),
    .Q_N(_01026_),
    .Q(net126));
 sg13g2_dfrbp_1 _16625_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net955),
    .D(\dp.ISRmux.d0[5] ),
    .Q_N(_01027_),
    .Q(net127));
 sg13g2_dfrbp_1 _16626_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net955),
    .D(\dp.ISRmux.d0[6] ),
    .Q_N(_01028_),
    .Q(net128));
 sg13g2_dfrbp_1 _16627_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net956),
    .D(\dp.ISRmux.d0[7] ),
    .Q_N(_01029_),
    .Q(net129));
 sg13g2_dfrbp_1 _16628_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net956),
    .D(\dp.ISRmux.d0[8] ),
    .Q_N(_01030_),
    .Q(net130));
 sg13g2_dfrbp_1 _16629_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net956),
    .D(\dp.ISRmux.d0[9] ),
    .Q_N(_01031_),
    .Q(net131));
 sg13g2_dfrbp_1 _16630_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net956),
    .D(\dp.ISRmux.d0[10] ),
    .Q_N(_01032_),
    .Q(net101));
 sg13g2_dfrbp_1 _16631_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net955),
    .D(\dp.ISRmux.d0[11] ),
    .Q_N(_01033_),
    .Q(net102));
 sg13g2_dfrbp_1 _16632_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net957),
    .D(\dp.ISRmux.d0[12] ),
    .Q_N(_01034_),
    .Q(net103));
 sg13g2_dfrbp_1 _16633_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net957),
    .D(\dp.ISRmux.d0[13] ),
    .Q_N(_01035_),
    .Q(net104));
 sg13g2_dfrbp_1 _16634_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net957),
    .D(\dp.ISRmux.d0[14] ),
    .Q_N(_01036_),
    .Q(net105));
 sg13g2_dfrbp_1 _16635_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net957),
    .D(\dp.ISRmux.d0[15] ),
    .Q_N(_01037_),
    .Q(net106));
 sg13g2_dfrbp_1 _16636_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net957),
    .D(\dp.ISRmux.d0[16] ),
    .Q_N(_01038_),
    .Q(net107));
 sg13g2_dfrbp_1 _16637_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net954),
    .D(\dp.ISRmux.d0[17] ),
    .Q_N(_01039_),
    .Q(net108));
 sg13g2_dfrbp_1 _16638_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net954),
    .D(\dp.ISRmux.d0[18] ),
    .Q_N(_01040_),
    .Q(net109));
 sg13g2_dfrbp_1 _16639_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net954),
    .D(\dp.ISRmux.d0[19] ),
    .Q_N(_01041_),
    .Q(net110));
 sg13g2_dfrbp_1 _16640_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net953),
    .D(\dp.ISRmux.d0[20] ),
    .Q_N(_01042_),
    .Q(net112));
 sg13g2_dfrbp_1 _16641_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net953),
    .D(\dp.ISRmux.d0[21] ),
    .Q_N(_01043_),
    .Q(net113));
 sg13g2_dfrbp_1 _16642_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net953),
    .D(\dp.ISRmux.d0[22] ),
    .Q_N(_01044_),
    .Q(net114));
 sg13g2_dfrbp_1 _16643_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net953),
    .D(\dp.ISRmux.d0[23] ),
    .Q_N(_01045_),
    .Q(net115));
 sg13g2_dfrbp_1 _16644_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net953),
    .D(\dp.ISRmux.d0[24] ),
    .Q_N(_01046_),
    .Q(net116));
 sg13g2_dfrbp_1 _16645_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net953),
    .D(\dp.ISRmux.d0[25] ),
    .Q_N(_01047_),
    .Q(net117));
 sg13g2_dfrbp_1 _16646_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net953),
    .D(\dp.ISRmux.d0[26] ),
    .Q_N(_01048_),
    .Q(net118));
 sg13g2_dfrbp_1 _16647_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net953),
    .D(\dp.ISRmux.d0[27] ),
    .Q_N(_01049_),
    .Q(net119));
 sg13g2_dfrbp_1 _16648_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net954),
    .D(\dp.ISRmux.d0[28] ),
    .Q_N(_01050_),
    .Q(net120));
 sg13g2_dfrbp_1 _16649_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net954),
    .D(\dp.ISRmux.d0[29] ),
    .Q_N(_01051_),
    .Q(net121));
 sg13g2_dfrbp_1 _16650_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net954),
    .D(\dp.ISRmux.d0[30] ),
    .Q_N(_01052_),
    .Q(net123));
 sg13g2_dfrbp_1 _16651_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net954),
    .D(\dp.ISRmux.d0[31] ),
    .Q_N(_08517_),
    .Q(net124));
 sg13g2_dfrbp_1 _16652_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01596_),
    .Q_N(_00009_),
    .Q(\dp.rf.rf[9][0] ));
 sg13g2_dfrbp_1 _16653_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_08518_),
    .D(_01597_),
    .Q_N(_00999_),
    .Q(\dp.rf.rf[9][1] ));
 sg13g2_dfrbp_1 _16654_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01598_),
    .Q_N(_00967_),
    .Q(\dp.rf.rf[9][2] ));
 sg13g2_dfrbp_1 _16655_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(_08518_),
    .D(_01599_),
    .Q_N(_00935_),
    .Q(\dp.rf.rf[9][3] ));
 sg13g2_dfrbp_1 _16656_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_08518_),
    .D(_01600_),
    .Q_N(_00903_),
    .Q(\dp.rf.rf[9][4] ));
 sg13g2_dfrbp_1 _16657_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_08518_),
    .D(_01601_),
    .Q_N(_00871_),
    .Q(\dp.rf.rf[9][5] ));
 sg13g2_dfrbp_1 _16658_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_08518_),
    .D(_01602_),
    .Q_N(_00839_),
    .Q(\dp.rf.rf[9][6] ));
 sg13g2_dfrbp_1 _16659_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01603_),
    .Q_N(_00807_),
    .Q(\dp.rf.rf[9][7] ));
 sg13g2_dfrbp_1 _16660_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(_08518_),
    .D(_01604_),
    .Q_N(_00775_),
    .Q(\dp.rf.rf[9][8] ));
 sg13g2_dfrbp_1 _16661_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01605_),
    .Q_N(_00743_),
    .Q(\dp.rf.rf[9][9] ));
 sg13g2_dfrbp_1 _16662_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01606_),
    .Q_N(_00711_),
    .Q(\dp.rf.rf[9][10] ));
 sg13g2_dfrbp_1 _16663_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01607_),
    .Q_N(_00679_),
    .Q(\dp.rf.rf[9][11] ));
 sg13g2_dfrbp_1 _16664_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01608_),
    .Q_N(_00647_),
    .Q(\dp.rf.rf[9][12] ));
 sg13g2_dfrbp_1 _16665_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_08518_),
    .D(_01609_),
    .Q_N(_00615_),
    .Q(\dp.rf.rf[9][13] ));
 sg13g2_dfrbp_1 _16666_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01610_),
    .Q_N(_00583_),
    .Q(\dp.rf.rf[9][14] ));
 sg13g2_dfrbp_1 _16667_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_08518_),
    .D(_01611_),
    .Q_N(_00551_),
    .Q(\dp.rf.rf[9][15] ));
 sg13g2_dfrbp_1 _16668_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_01612_),
    .Q_N(_00519_),
    .Q(\dp.rf.rf[9][16] ));
 sg13g2_dfrbp_1 _16669_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(_08518_),
    .D(_01613_),
    .Q_N(_00487_),
    .Q(\dp.rf.rf[9][17] ));
 sg13g2_dfrbp_1 _16670_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(_01614_),
    .Q_N(_00456_),
    .Q(\dp.rf.rf[9][18] ));
 sg13g2_dfrbp_1 _16671_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(_01615_),
    .Q_N(_00424_),
    .Q(\dp.rf.rf[9][19] ));
 sg13g2_dfrbp_1 _16672_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(_08518_),
    .D(_01616_),
    .Q_N(_00393_),
    .Q(\dp.rf.rf[9][20] ));
 sg13g2_dfrbp_1 _16673_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01617_),
    .Q_N(_00361_),
    .Q(\dp.rf.rf[9][21] ));
 sg13g2_dfrbp_1 _16674_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01618_),
    .Q_N(_00329_),
    .Q(\dp.rf.rf[9][22] ));
 sg13g2_dfrbp_1 _16675_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01619_),
    .Q_N(_00297_),
    .Q(\dp.rf.rf[9][23] ));
 sg13g2_dfrbp_1 _16676_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01620_),
    .Q_N(_00265_),
    .Q(\dp.rf.rf[9][24] ));
 sg13g2_dfrbp_1 _16677_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01621_),
    .Q_N(_00233_),
    .Q(\dp.rf.rf[9][25] ));
 sg13g2_dfrbp_1 _16678_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_01622_),
    .Q_N(_00201_),
    .Q(\dp.rf.rf[9][26] ));
 sg13g2_dfrbp_1 _16679_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_01623_),
    .Q_N(_00169_),
    .Q(\dp.rf.rf[9][27] ));
 sg13g2_dfrbp_1 _16680_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01624_),
    .Q_N(_00137_),
    .Q(\dp.rf.rf[9][28] ));
 sg13g2_dfrbp_1 _16681_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01625_),
    .Q_N(_00105_),
    .Q(\dp.rf.rf[9][29] ));
 sg13g2_dfrbp_1 _16682_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_01626_),
    .Q_N(_00073_),
    .Q(\dp.rf.rf[9][30] ));
 sg13g2_dfrbp_1 _16683_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_01627_),
    .Q_N(_00041_),
    .Q(\dp.rf.rf[9][31] ));
 sg13g2_dfrbp_1 _16684_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_08518_),
    .D(_01628_),
    .Q_N(_00022_),
    .Q(\dp.rf.rf[22][0] ));
 sg13g2_dfrbp_1 _16685_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01629_),
    .Q_N(_01012_),
    .Q(\dp.rf.rf[22][1] ));
 sg13g2_dfrbp_1 _16686_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01630_),
    .Q_N(_00980_),
    .Q(\dp.rf.rf[22][2] ));
 sg13g2_dfrbp_1 _16687_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01631_),
    .Q_N(_00948_),
    .Q(\dp.rf.rf[22][3] ));
 sg13g2_dfrbp_1 _16688_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(_01632_),
    .Q_N(_00916_),
    .Q(\dp.rf.rf[22][4] ));
 sg13g2_dfrbp_1 _16689_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_08518_),
    .D(_01633_),
    .Q_N(_00884_),
    .Q(\dp.rf.rf[22][5] ));
 sg13g2_dfrbp_1 _16690_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01634_),
    .Q_N(_00852_),
    .Q(\dp.rf.rf[22][6] ));
 sg13g2_dfrbp_1 _16691_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01635_),
    .Q_N(_00820_),
    .Q(\dp.rf.rf[22][7] ));
 sg13g2_dfrbp_1 _16692_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01636_),
    .Q_N(_00788_),
    .Q(\dp.rf.rf[22][8] ));
 sg13g2_dfrbp_1 _16693_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01637_),
    .Q_N(_00756_),
    .Q(\dp.rf.rf[22][9] ));
 sg13g2_dfrbp_1 _16694_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01638_),
    .Q_N(_00724_),
    .Q(\dp.rf.rf[22][10] ));
 sg13g2_dfrbp_1 _16695_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_01639_),
    .Q_N(_00692_),
    .Q(\dp.rf.rf[22][11] ));
 sg13g2_dfrbp_1 _16696_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_08518_),
    .D(_01640_),
    .Q_N(_00660_),
    .Q(\dp.rf.rf[22][12] ));
 sg13g2_dfrbp_1 _16697_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_08518_),
    .D(_01641_),
    .Q_N(_00628_),
    .Q(\dp.rf.rf[22][13] ));
 sg13g2_dfrbp_1 _16698_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01642_),
    .Q_N(_00596_),
    .Q(\dp.rf.rf[22][14] ));
 sg13g2_dfrbp_1 _16699_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01643_),
    .Q_N(_00564_),
    .Q(\dp.rf.rf[22][15] ));
 sg13g2_dfrbp_1 _16700_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01644_),
    .Q_N(_00532_),
    .Q(\dp.rf.rf[22][16] ));
 sg13g2_dfrbp_1 _16701_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(_08518_),
    .D(_01645_),
    .Q_N(_00500_),
    .Q(\dp.rf.rf[22][17] ));
 sg13g2_dfrbp_1 _16702_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_01646_),
    .Q_N(_00469_),
    .Q(\dp.rf.rf[22][18] ));
 sg13g2_dfrbp_1 _16703_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01647_),
    .Q_N(_00437_),
    .Q(\dp.rf.rf[22][19] ));
 sg13g2_dfrbp_1 _16704_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(_08518_),
    .D(_01648_),
    .Q_N(_00406_),
    .Q(\dp.rf.rf[22][20] ));
 sg13g2_dfrbp_1 _16705_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01649_),
    .Q_N(_00374_),
    .Q(\dp.rf.rf[22][21] ));
 sg13g2_dfrbp_1 _16706_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01650_),
    .Q_N(_00342_),
    .Q(\dp.rf.rf[22][22] ));
 sg13g2_dfrbp_1 _16707_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01651_),
    .Q_N(_00310_),
    .Q(\dp.rf.rf[22][23] ));
 sg13g2_dfrbp_1 _16708_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(_08518_),
    .D(_01652_),
    .Q_N(_00278_),
    .Q(\dp.rf.rf[22][24] ));
 sg13g2_dfrbp_1 _16709_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01653_),
    .Q_N(_00246_),
    .Q(\dp.rf.rf[22][25] ));
 sg13g2_dfrbp_1 _16710_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01654_),
    .Q_N(_00214_),
    .Q(\dp.rf.rf[22][26] ));
 sg13g2_dfrbp_1 _16711_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01655_),
    .Q_N(_00182_),
    .Q(\dp.rf.rf[22][27] ));
 sg13g2_dfrbp_1 _16712_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01656_),
    .Q_N(_00150_),
    .Q(\dp.rf.rf[22][28] ));
 sg13g2_dfrbp_1 _16713_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01657_),
    .Q_N(_00118_),
    .Q(\dp.rf.rf[22][29] ));
 sg13g2_dfrbp_1 _16714_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01658_),
    .Q_N(_00086_),
    .Q(\dp.rf.rf[22][30] ));
 sg13g2_dfrbp_1 _16715_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01659_),
    .Q_N(_00054_),
    .Q(\dp.rf.rf[22][31] ));
 sg13g2_dfrbp_1 _16716_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_08518_),
    .D(_01660_),
    .Q_N(_00025_),
    .Q(\dp.rf.rf[25][0] ));
 sg13g2_dfrbp_1 _16717_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01661_),
    .Q_N(_01015_),
    .Q(\dp.rf.rf[25][1] ));
 sg13g2_dfrbp_1 _16718_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01662_),
    .Q_N(_00983_),
    .Q(\dp.rf.rf[25][2] ));
 sg13g2_dfrbp_1 _16719_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01663_),
    .Q_N(_00951_),
    .Q(\dp.rf.rf[25][3] ));
 sg13g2_dfrbp_1 _16720_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01664_),
    .Q_N(_00919_),
    .Q(\dp.rf.rf[25][4] ));
 sg13g2_dfrbp_1 _16721_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01665_),
    .Q_N(_00887_),
    .Q(\dp.rf.rf[25][5] ));
 sg13g2_dfrbp_1 _16722_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01666_),
    .Q_N(_00855_),
    .Q(\dp.rf.rf[25][6] ));
 sg13g2_dfrbp_1 _16723_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01667_),
    .Q_N(_00823_),
    .Q(\dp.rf.rf[25][7] ));
 sg13g2_dfrbp_1 _16724_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01668_),
    .Q_N(_00791_),
    .Q(\dp.rf.rf[25][8] ));
 sg13g2_dfrbp_1 _16725_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01669_),
    .Q_N(_00759_),
    .Q(\dp.rf.rf[25][9] ));
 sg13g2_dfrbp_1 _16726_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01670_),
    .Q_N(_00727_),
    .Q(\dp.rf.rf[25][10] ));
 sg13g2_dfrbp_1 _16727_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01671_),
    .Q_N(_00695_),
    .Q(\dp.rf.rf[25][11] ));
 sg13g2_dfrbp_1 _16728_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_08518_),
    .D(_01672_),
    .Q_N(_00663_),
    .Q(\dp.rf.rf[25][12] ));
 sg13g2_dfrbp_1 _16729_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(_08518_),
    .D(_01673_),
    .Q_N(_00631_),
    .Q(\dp.rf.rf[25][13] ));
 sg13g2_dfrbp_1 _16730_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(_08518_),
    .D(_01674_),
    .Q_N(_00599_),
    .Q(\dp.rf.rf[25][14] ));
 sg13g2_dfrbp_1 _16731_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_08518_),
    .D(_01675_),
    .Q_N(_00567_),
    .Q(\dp.rf.rf[25][15] ));
 sg13g2_dfrbp_1 _16732_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01676_),
    .Q_N(_00535_),
    .Q(\dp.rf.rf[25][16] ));
 sg13g2_dfrbp_1 _16733_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(_08518_),
    .D(_01677_),
    .Q_N(_00503_),
    .Q(\dp.rf.rf[25][17] ));
 sg13g2_dfrbp_1 _16734_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01678_),
    .Q_N(_00472_),
    .Q(\dp.rf.rf[25][18] ));
 sg13g2_dfrbp_1 _16735_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(_01679_),
    .Q_N(_00440_),
    .Q(\dp.rf.rf[25][19] ));
 sg13g2_dfrbp_1 _16736_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01680_),
    .Q_N(_00409_),
    .Q(\dp.rf.rf[25][20] ));
 sg13g2_dfrbp_1 _16737_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01681_),
    .Q_N(_00377_),
    .Q(\dp.rf.rf[25][21] ));
 sg13g2_dfrbp_1 _16738_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(_08518_),
    .D(_01682_),
    .Q_N(_00345_),
    .Q(\dp.rf.rf[25][22] ));
 sg13g2_dfrbp_1 _16739_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_01683_),
    .Q_N(_00313_),
    .Q(\dp.rf.rf[25][23] ));
 sg13g2_dfrbp_1 _16740_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(_08518_),
    .D(_01684_),
    .Q_N(_00281_),
    .Q(\dp.rf.rf[25][24] ));
 sg13g2_dfrbp_1 _16741_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_01685_),
    .Q_N(_00249_),
    .Q(\dp.rf.rf[25][25] ));
 sg13g2_dfrbp_1 _16742_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01686_),
    .Q_N(_00217_),
    .Q(\dp.rf.rf[25][26] ));
 sg13g2_dfrbp_1 _16743_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01687_),
    .Q_N(_00185_),
    .Q(\dp.rf.rf[25][27] ));
 sg13g2_dfrbp_1 _16744_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01688_),
    .Q_N(_00153_),
    .Q(\dp.rf.rf[25][28] ));
 sg13g2_dfrbp_1 _16745_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01689_),
    .Q_N(_00121_),
    .Q(\dp.rf.rf[25][29] ));
 sg13g2_dfrbp_1 _16746_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01690_),
    .Q_N(_00089_),
    .Q(\dp.rf.rf[25][30] ));
 sg13g2_dfrbp_1 _16747_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01691_),
    .Q_N(_00057_),
    .Q(\dp.rf.rf[25][31] ));
 sg13g2_dfrbp_1 _16748_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_08518_),
    .D(_01692_),
    .Q_N(_00026_),
    .Q(\dp.rf.rf[26][0] ));
 sg13g2_dfrbp_1 _16749_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01693_),
    .Q_N(_01016_),
    .Q(\dp.rf.rf[26][1] ));
 sg13g2_dfrbp_1 _16750_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01694_),
    .Q_N(_00984_),
    .Q(\dp.rf.rf[26][2] ));
 sg13g2_dfrbp_1 _16751_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01695_),
    .Q_N(_00952_),
    .Q(\dp.rf.rf[26][3] ));
 sg13g2_dfrbp_1 _16752_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01696_),
    .Q_N(_00920_),
    .Q(\dp.rf.rf[26][4] ));
 sg13g2_dfrbp_1 _16753_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01697_),
    .Q_N(_00888_),
    .Q(\dp.rf.rf[26][5] ));
 sg13g2_dfrbp_1 _16754_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01698_),
    .Q_N(_00856_),
    .Q(\dp.rf.rf[26][6] ));
 sg13g2_dfrbp_1 _16755_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01699_),
    .Q_N(_00824_),
    .Q(\dp.rf.rf[26][7] ));
 sg13g2_dfrbp_1 _16756_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01700_),
    .Q_N(_00792_),
    .Q(\dp.rf.rf[26][8] ));
 sg13g2_dfrbp_1 _16757_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01701_),
    .Q_N(_00760_),
    .Q(\dp.rf.rf[26][9] ));
 sg13g2_dfrbp_1 _16758_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01702_),
    .Q_N(_00728_),
    .Q(\dp.rf.rf[26][10] ));
 sg13g2_dfrbp_1 _16759_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01703_),
    .Q_N(_00696_),
    .Q(\dp.rf.rf[26][11] ));
 sg13g2_dfrbp_1 _16760_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_08518_),
    .D(_01704_),
    .Q_N(_00664_),
    .Q(\dp.rf.rf[26][12] ));
 sg13g2_dfrbp_1 _16761_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(_08518_),
    .D(_01705_),
    .Q_N(_00632_),
    .Q(\dp.rf.rf[26][13] ));
 sg13g2_dfrbp_1 _16762_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(_08518_),
    .D(_01706_),
    .Q_N(_00600_),
    .Q(\dp.rf.rf[26][14] ));
 sg13g2_dfrbp_1 _16763_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01707_),
    .Q_N(_00568_),
    .Q(\dp.rf.rf[26][15] ));
 sg13g2_dfrbp_1 _16764_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01708_),
    .Q_N(_00536_),
    .Q(\dp.rf.rf[26][16] ));
 sg13g2_dfrbp_1 _16765_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(_08518_),
    .D(_01709_),
    .Q_N(_00504_),
    .Q(\dp.rf.rf[26][17] ));
 sg13g2_dfrbp_1 _16766_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_01710_),
    .Q_N(_00473_),
    .Q(\dp.rf.rf[26][18] ));
 sg13g2_dfrbp_1 _16767_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(_01711_),
    .Q_N(_00441_),
    .Q(\dp.rf.rf[26][19] ));
 sg13g2_dfrbp_1 _16768_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01712_),
    .Q_N(_00410_),
    .Q(\dp.rf.rf[26][20] ));
 sg13g2_dfrbp_1 _16769_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01713_),
    .Q_N(_00378_),
    .Q(\dp.rf.rf[26][21] ));
 sg13g2_dfrbp_1 _16770_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01714_),
    .Q_N(_00346_),
    .Q(\dp.rf.rf[26][22] ));
 sg13g2_dfrbp_1 _16771_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_01715_),
    .Q_N(_00314_),
    .Q(\dp.rf.rf[26][23] ));
 sg13g2_dfrbp_1 _16772_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(_08518_),
    .D(_01716_),
    .Q_N(_00282_),
    .Q(\dp.rf.rf[26][24] ));
 sg13g2_dfrbp_1 _16773_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_01717_),
    .Q_N(_00250_),
    .Q(\dp.rf.rf[26][25] ));
 sg13g2_dfrbp_1 _16774_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01718_),
    .Q_N(_00218_),
    .Q(\dp.rf.rf[26][26] ));
 sg13g2_dfrbp_1 _16775_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01719_),
    .Q_N(_00186_),
    .Q(\dp.rf.rf[26][27] ));
 sg13g2_dfrbp_1 _16776_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01720_),
    .Q_N(_00154_),
    .Q(\dp.rf.rf[26][28] ));
 sg13g2_dfrbp_1 _16777_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01721_),
    .Q_N(_00122_),
    .Q(\dp.rf.rf[26][29] ));
 sg13g2_dfrbp_1 _16778_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01722_),
    .Q_N(_00090_),
    .Q(\dp.rf.rf[26][30] ));
 sg13g2_dfrbp_1 _16779_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01723_),
    .Q_N(_00058_),
    .Q(\dp.rf.rf[26][31] ));
 sg13g2_dfrbp_1 _16780_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_01724_),
    .Q_N(_00028_),
    .Q(\dp.rf.rf[28][0] ));
 sg13g2_dfrbp_1 _16781_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01725_),
    .Q_N(_01018_),
    .Q(\dp.rf.rf[28][1] ));
 sg13g2_dfrbp_1 _16782_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01726_),
    .Q_N(_00986_),
    .Q(\dp.rf.rf[28][2] ));
 sg13g2_dfrbp_1 _16783_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01727_),
    .Q_N(_00954_),
    .Q(\dp.rf.rf[28][3] ));
 sg13g2_dfrbp_1 _16784_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01728_),
    .Q_N(_00922_),
    .Q(\dp.rf.rf[28][4] ));
 sg13g2_dfrbp_1 _16785_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01729_),
    .Q_N(_00890_),
    .Q(\dp.rf.rf[28][5] ));
 sg13g2_dfrbp_1 _16786_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01730_),
    .Q_N(_00858_),
    .Q(\dp.rf.rf[28][6] ));
 sg13g2_dfrbp_1 _16787_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01731_),
    .Q_N(_00826_),
    .Q(\dp.rf.rf[28][7] ));
 sg13g2_dfrbp_1 _16788_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01732_),
    .Q_N(_00794_),
    .Q(\dp.rf.rf[28][8] ));
 sg13g2_dfrbp_1 _16789_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_08518_),
    .D(_01733_),
    .Q_N(_00762_),
    .Q(\dp.rf.rf[28][9] ));
 sg13g2_dfrbp_1 _16790_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01734_),
    .Q_N(_00730_),
    .Q(\dp.rf.rf[28][10] ));
 sg13g2_dfrbp_1 _16791_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01735_),
    .Q_N(_00698_),
    .Q(\dp.rf.rf[28][11] ));
 sg13g2_dfrbp_1 _16792_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_08518_),
    .D(_01736_),
    .Q_N(_00666_),
    .Q(\dp.rf.rf[28][12] ));
 sg13g2_dfrbp_1 _16793_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(_08518_),
    .D(_01737_),
    .Q_N(_00634_),
    .Q(\dp.rf.rf[28][13] ));
 sg13g2_dfrbp_1 _16794_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(_01738_),
    .Q_N(_00602_),
    .Q(\dp.rf.rf[28][14] ));
 sg13g2_dfrbp_1 _16795_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_08518_),
    .D(_01739_),
    .Q_N(_00570_),
    .Q(\dp.rf.rf[28][15] ));
 sg13g2_dfrbp_1 _16796_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01740_),
    .Q_N(_00538_),
    .Q(\dp.rf.rf[28][16] ));
 sg13g2_dfrbp_1 _16797_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(_08518_),
    .D(_01741_),
    .Q_N(_00506_),
    .Q(\dp.rf.rf[28][17] ));
 sg13g2_dfrbp_1 _16798_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01742_),
    .Q_N(_00475_),
    .Q(\dp.rf.rf[28][18] ));
 sg13g2_dfrbp_1 _16799_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_08518_),
    .D(_01743_),
    .Q_N(_00443_),
    .Q(\dp.rf.rf[28][19] ));
 sg13g2_dfrbp_1 _16800_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(_08518_),
    .D(_01744_),
    .Q_N(_00412_),
    .Q(\dp.rf.rf[28][20] ));
 sg13g2_dfrbp_1 _16801_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01745_),
    .Q_N(_00380_),
    .Q(\dp.rf.rf[28][21] ));
 sg13g2_dfrbp_1 _16802_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01746_),
    .Q_N(_00348_),
    .Q(\dp.rf.rf[28][22] ));
 sg13g2_dfrbp_1 _16803_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01747_),
    .Q_N(_00316_),
    .Q(\dp.rf.rf[28][23] ));
 sg13g2_dfrbp_1 _16804_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01748_),
    .Q_N(_00284_),
    .Q(\dp.rf.rf[28][24] ));
 sg13g2_dfrbp_1 _16805_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01749_),
    .Q_N(_00252_),
    .Q(\dp.rf.rf[28][25] ));
 sg13g2_dfrbp_1 _16806_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(_08518_),
    .D(_01750_),
    .Q_N(_00220_),
    .Q(\dp.rf.rf[28][26] ));
 sg13g2_dfrbp_1 _16807_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(_08518_),
    .D(_01751_),
    .Q_N(_00188_),
    .Q(\dp.rf.rf[28][27] ));
 sg13g2_dfrbp_1 _16808_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_01752_),
    .Q_N(_00156_),
    .Q(\dp.rf.rf[28][28] ));
 sg13g2_dfrbp_1 _16809_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(_08518_),
    .D(_01753_),
    .Q_N(_00124_),
    .Q(\dp.rf.rf[28][29] ));
 sg13g2_dfrbp_1 _16810_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(_08518_),
    .D(_01754_),
    .Q_N(_00092_),
    .Q(\dp.rf.rf[28][30] ));
 sg13g2_dfrbp_1 _16811_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01755_),
    .Q_N(_00060_),
    .Q(\dp.rf.rf[28][31] ));
 sg13g2_dfrbp_1 _16812_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_08518_),
    .D(_01756_),
    .Q_N(_00027_),
    .Q(\dp.rf.rf[27][0] ));
 sg13g2_dfrbp_1 _16813_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01757_),
    .Q_N(_01017_),
    .Q(\dp.rf.rf[27][1] ));
 sg13g2_dfrbp_1 _16814_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01758_),
    .Q_N(_00985_),
    .Q(\dp.rf.rf[27][2] ));
 sg13g2_dfrbp_1 _16815_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01759_),
    .Q_N(_00953_),
    .Q(\dp.rf.rf[27][3] ));
 sg13g2_dfrbp_1 _16816_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01760_),
    .Q_N(_00921_),
    .Q(\dp.rf.rf[27][4] ));
 sg13g2_dfrbp_1 _16817_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_08518_),
    .D(_01761_),
    .Q_N(_00889_),
    .Q(\dp.rf.rf[27][5] ));
 sg13g2_dfrbp_1 _16818_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01762_),
    .Q_N(_00857_),
    .Q(\dp.rf.rf[27][6] ));
 sg13g2_dfrbp_1 _16819_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01763_),
    .Q_N(_00825_),
    .Q(\dp.rf.rf[27][7] ));
 sg13g2_dfrbp_1 _16820_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01764_),
    .Q_N(_00793_),
    .Q(\dp.rf.rf[27][8] ));
 sg13g2_dfrbp_1 _16821_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01765_),
    .Q_N(_00761_),
    .Q(\dp.rf.rf[27][9] ));
 sg13g2_dfrbp_1 _16822_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01766_),
    .Q_N(_00729_),
    .Q(\dp.rf.rf[27][10] ));
 sg13g2_dfrbp_1 _16823_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01767_),
    .Q_N(_00697_),
    .Q(\dp.rf.rf[27][11] ));
 sg13g2_dfrbp_1 _16824_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_08518_),
    .D(_01768_),
    .Q_N(_00665_),
    .Q(\dp.rf.rf[27][12] ));
 sg13g2_dfrbp_1 _16825_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(_08518_),
    .D(_01769_),
    .Q_N(_00633_),
    .Q(\dp.rf.rf[27][13] ));
 sg13g2_dfrbp_1 _16826_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(_08518_),
    .D(_01770_),
    .Q_N(_00601_),
    .Q(\dp.rf.rf[27][14] ));
 sg13g2_dfrbp_1 _16827_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_08518_),
    .D(_01771_),
    .Q_N(_00569_),
    .Q(\dp.rf.rf[27][15] ));
 sg13g2_dfrbp_1 _16828_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01772_),
    .Q_N(_00537_),
    .Q(\dp.rf.rf[27][16] ));
 sg13g2_dfrbp_1 _16829_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(_08518_),
    .D(_01773_),
    .Q_N(_00505_),
    .Q(\dp.rf.rf[27][17] ));
 sg13g2_dfrbp_1 _16830_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01774_),
    .Q_N(_00474_),
    .Q(\dp.rf.rf[27][18] ));
 sg13g2_dfrbp_1 _16831_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_08518_),
    .D(_01775_),
    .Q_N(_00442_),
    .Q(\dp.rf.rf[27][19] ));
 sg13g2_dfrbp_1 _16832_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01776_),
    .Q_N(_00411_),
    .Q(\dp.rf.rf[27][20] ));
 sg13g2_dfrbp_1 _16833_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01777_),
    .Q_N(_00379_),
    .Q(\dp.rf.rf[27][21] ));
 sg13g2_dfrbp_1 _16834_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(_08518_),
    .D(_01778_),
    .Q_N(_00347_),
    .Q(\dp.rf.rf[27][22] ));
 sg13g2_dfrbp_1 _16835_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_01779_),
    .Q_N(_00315_),
    .Q(\dp.rf.rf[27][23] ));
 sg13g2_dfrbp_1 _16836_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(_08518_),
    .D(_01780_),
    .Q_N(_00283_),
    .Q(\dp.rf.rf[27][24] ));
 sg13g2_dfrbp_1 _16837_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_01781_),
    .Q_N(_00251_),
    .Q(\dp.rf.rf[27][25] ));
 sg13g2_dfrbp_1 _16838_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01782_),
    .Q_N(_00219_),
    .Q(\dp.rf.rf[27][26] ));
 sg13g2_dfrbp_1 _16839_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01783_),
    .Q_N(_00187_),
    .Q(\dp.rf.rf[27][27] ));
 sg13g2_dfrbp_1 _16840_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01784_),
    .Q_N(_00155_),
    .Q(\dp.rf.rf[27][28] ));
 sg13g2_dfrbp_1 _16841_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01785_),
    .Q_N(_00123_),
    .Q(\dp.rf.rf[27][29] ));
 sg13g2_dfrbp_1 _16842_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01786_),
    .Q_N(_00091_),
    .Q(\dp.rf.rf[27][30] ));
 sg13g2_dfrbp_1 _16843_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01787_),
    .Q_N(_00059_),
    .Q(\dp.rf.rf[27][31] ));
 sg13g2_dfrbp_1 _16844_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_08518_),
    .D(_01788_),
    .Q_N(_00002_),
    .Q(\dp.rf.rf[2][0] ));
 sg13g2_dfrbp_1 _16845_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01789_),
    .Q_N(_00992_),
    .Q(\dp.rf.rf[2][1] ));
 sg13g2_dfrbp_1 _16846_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01790_),
    .Q_N(_00960_),
    .Q(\dp.rf.rf[2][2] ));
 sg13g2_dfrbp_1 _16847_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_01791_),
    .Q_N(_00928_),
    .Q(\dp.rf.rf[2][3] ));
 sg13g2_dfrbp_1 _16848_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_08518_),
    .D(_01792_),
    .Q_N(_00896_),
    .Q(\dp.rf.rf[2][4] ));
 sg13g2_dfrbp_1 _16849_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_08518_),
    .D(_01793_),
    .Q_N(_00864_),
    .Q(\dp.rf.rf[2][5] ));
 sg13g2_dfrbp_1 _16850_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01794_),
    .Q_N(_00832_),
    .Q(\dp.rf.rf[2][6] ));
 sg13g2_dfrbp_1 _16851_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01795_),
    .Q_N(_00800_),
    .Q(\dp.rf.rf[2][7] ));
 sg13g2_dfrbp_1 _16852_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_01796_),
    .Q_N(_00768_),
    .Q(\dp.rf.rf[2][8] ));
 sg13g2_dfrbp_1 _16853_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_01797_),
    .Q_N(_00736_),
    .Q(\dp.rf.rf[2][9] ));
 sg13g2_dfrbp_1 _16854_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01798_),
    .Q_N(_00704_),
    .Q(\dp.rf.rf[2][10] ));
 sg13g2_dfrbp_1 _16855_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01799_),
    .Q_N(_00672_),
    .Q(\dp.rf.rf[2][11] ));
 sg13g2_dfrbp_1 _16856_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_01800_),
    .Q_N(_00640_),
    .Q(\dp.rf.rf[2][12] ));
 sg13g2_dfrbp_1 _16857_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_08518_),
    .D(_01801_),
    .Q_N(_00608_),
    .Q(\dp.rf.rf[2][13] ));
 sg13g2_dfrbp_1 _16858_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01802_),
    .Q_N(_00576_),
    .Q(\dp.rf.rf[2][14] ));
 sg13g2_dfrbp_1 _16859_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_01803_),
    .Q_N(_00544_),
    .Q(\dp.rf.rf[2][15] ));
 sg13g2_dfrbp_1 _16860_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_01804_),
    .Q_N(_00512_),
    .Q(\dp.rf.rf[2][16] ));
 sg13g2_dfrbp_1 _16861_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(_08518_),
    .D(_01805_),
    .Q_N(_00480_),
    .Q(\dp.rf.rf[2][17] ));
 sg13g2_dfrbp_1 _16862_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(_01806_),
    .Q_N(_00449_),
    .Q(\dp.rf.rf[2][18] ));
 sg13g2_dfrbp_1 _16863_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_08518_),
    .D(_01807_),
    .Q_N(_00417_),
    .Q(\dp.rf.rf[2][19] ));
 sg13g2_dfrbp_1 _16864_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(_08518_),
    .D(_01808_),
    .Q_N(_00386_),
    .Q(\dp.rf.rf[2][20] ));
 sg13g2_dfrbp_1 _16865_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_01809_),
    .Q_N(_00354_),
    .Q(\dp.rf.rf[2][21] ));
 sg13g2_dfrbp_1 _16866_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01810_),
    .Q_N(_00322_),
    .Q(\dp.rf.rf[2][22] ));
 sg13g2_dfrbp_1 _16867_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_08518_),
    .D(_01811_),
    .Q_N(_00290_),
    .Q(\dp.rf.rf[2][23] ));
 sg13g2_dfrbp_1 _16868_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(_08518_),
    .D(_01812_),
    .Q_N(_00258_),
    .Q(\dp.rf.rf[2][24] ));
 sg13g2_dfrbp_1 _16869_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_01813_),
    .Q_N(_00226_),
    .Q(\dp.rf.rf[2][25] ));
 sg13g2_dfrbp_1 _16870_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(_08518_),
    .D(_01814_),
    .Q_N(_00194_),
    .Q(\dp.rf.rf[2][26] ));
 sg13g2_dfrbp_1 _16871_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01815_),
    .Q_N(_00162_),
    .Q(\dp.rf.rf[2][27] ));
 sg13g2_dfrbp_1 _16872_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_01816_),
    .Q_N(_00130_),
    .Q(\dp.rf.rf[2][28] ));
 sg13g2_dfrbp_1 _16873_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(_08518_),
    .D(_01817_),
    .Q_N(_00098_),
    .Q(\dp.rf.rf[2][29] ));
 sg13g2_dfrbp_1 _16874_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01818_),
    .Q_N(_00066_),
    .Q(\dp.rf.rf[2][30] ));
 sg13g2_dfrbp_1 _16875_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_08518_),
    .D(_01819_),
    .Q_N(_00034_),
    .Q(\dp.rf.rf[2][31] ));
 sg13g2_dfrbp_1 _16876_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_08518_),
    .D(_01820_),
    .Q_N(_00030_),
    .Q(\dp.rf.rf[30][0] ));
 sg13g2_dfrbp_1 _16877_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01821_),
    .Q_N(_01020_),
    .Q(\dp.rf.rf[30][1] ));
 sg13g2_dfrbp_1 _16878_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01822_),
    .Q_N(_00988_),
    .Q(\dp.rf.rf[30][2] ));
 sg13g2_dfrbp_1 _16879_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(_08518_),
    .D(_01823_),
    .Q_N(_00956_),
    .Q(\dp.rf.rf[30][3] ));
 sg13g2_dfrbp_1 _16880_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(_08518_),
    .D(_01824_),
    .Q_N(_00924_),
    .Q(\dp.rf.rf[30][4] ));
 sg13g2_dfrbp_1 _16881_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01825_),
    .Q_N(_00892_),
    .Q(\dp.rf.rf[30][5] ));
 sg13g2_dfrbp_1 _16882_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01826_),
    .Q_N(_00860_),
    .Q(\dp.rf.rf[30][6] ));
 sg13g2_dfrbp_1 _16883_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01827_),
    .Q_N(_00828_),
    .Q(\dp.rf.rf[30][7] ));
 sg13g2_dfrbp_1 _16884_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01828_),
    .Q_N(_00796_),
    .Q(\dp.rf.rf[30][8] ));
 sg13g2_dfrbp_1 _16885_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01829_),
    .Q_N(_00764_),
    .Q(\dp.rf.rf[30][9] ));
 sg13g2_dfrbp_1 _16886_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_08518_),
    .D(_01830_),
    .Q_N(_00732_),
    .Q(\dp.rf.rf[30][10] ));
 sg13g2_dfrbp_1 _16887_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01831_),
    .Q_N(_00700_),
    .Q(\dp.rf.rf[30][11] ));
 sg13g2_dfrbp_1 _16888_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_08518_),
    .D(_01832_),
    .Q_N(_00668_),
    .Q(\dp.rf.rf[30][12] ));
 sg13g2_dfrbp_1 _16889_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(_08518_),
    .D(_01833_),
    .Q_N(_00636_),
    .Q(\dp.rf.rf[30][13] ));
 sg13g2_dfrbp_1 _16890_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01834_),
    .Q_N(_00604_),
    .Q(\dp.rf.rf[30][14] ));
 sg13g2_dfrbp_1 _16891_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(_08518_),
    .D(_01835_),
    .Q_N(_00572_),
    .Q(\dp.rf.rf[30][15] ));
 sg13g2_dfrbp_1 _16892_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_08518_),
    .D(_01836_),
    .Q_N(_00540_),
    .Q(\dp.rf.rf[30][16] ));
 sg13g2_dfrbp_1 _16893_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(_08518_),
    .D(_01837_),
    .Q_N(_00508_),
    .Q(\dp.rf.rf[30][17] ));
 sg13g2_dfrbp_1 _16894_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01838_),
    .Q_N(_00477_),
    .Q(\dp.rf.rf[30][18] ));
 sg13g2_dfrbp_1 _16895_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01839_),
    .Q_N(_00445_),
    .Q(\dp.rf.rf[30][19] ));
 sg13g2_dfrbp_1 _16896_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(_08518_),
    .D(_01840_),
    .Q_N(_00414_),
    .Q(\dp.rf.rf[30][20] ));
 sg13g2_dfrbp_1 _16897_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01841_),
    .Q_N(_00382_),
    .Q(\dp.rf.rf[30][21] ));
 sg13g2_dfrbp_1 _16898_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01842_),
    .Q_N(_00350_),
    .Q(\dp.rf.rf[30][22] ));
 sg13g2_dfrbp_1 _16899_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01843_),
    .Q_N(_00318_),
    .Q(\dp.rf.rf[30][23] ));
 sg13g2_dfrbp_1 _16900_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(_08518_),
    .D(_01844_),
    .Q_N(_00286_),
    .Q(\dp.rf.rf[30][24] ));
 sg13g2_dfrbp_1 _16901_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01845_),
    .Q_N(_00254_),
    .Q(\dp.rf.rf[30][25] ));
 sg13g2_dfrbp_1 _16902_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01846_),
    .Q_N(_00222_),
    .Q(\dp.rf.rf[30][26] ));
 sg13g2_dfrbp_1 _16903_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01847_),
    .Q_N(_00190_),
    .Q(\dp.rf.rf[30][27] ));
 sg13g2_dfrbp_1 _16904_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_01848_),
    .Q_N(_00158_),
    .Q(\dp.rf.rf[30][28] ));
 sg13g2_dfrbp_1 _16905_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01849_),
    .Q_N(_00126_),
    .Q(\dp.rf.rf[30][29] ));
 sg13g2_dfrbp_1 _16906_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(_08518_),
    .D(_01850_),
    .Q_N(_00094_),
    .Q(\dp.rf.rf[30][30] ));
 sg13g2_dfrbp_1 _16907_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01851_),
    .Q_N(_00062_),
    .Q(\dp.rf.rf[30][31] ));
 sg13g2_dfrbp_1 _16908_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(_08518_),
    .D(_01852_),
    .Q_N(_00024_),
    .Q(\dp.rf.rf[24][0] ));
 sg13g2_dfrbp_1 _16909_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01853_),
    .Q_N(_01014_),
    .Q(\dp.rf.rf[24][1] ));
 sg13g2_dfrbp_1 _16910_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01854_),
    .Q_N(_00982_),
    .Q(\dp.rf.rf[24][2] ));
 sg13g2_dfrbp_1 _16911_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01855_),
    .Q_N(_00950_),
    .Q(\dp.rf.rf[24][3] ));
 sg13g2_dfrbp_1 _16912_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01856_),
    .Q_N(_00918_),
    .Q(\dp.rf.rf[24][4] ));
 sg13g2_dfrbp_1 _16913_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(_08518_),
    .D(_01857_),
    .Q_N(_00886_),
    .Q(\dp.rf.rf[24][5] ));
 sg13g2_dfrbp_1 _16914_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01858_),
    .Q_N(_00854_),
    .Q(\dp.rf.rf[24][6] ));
 sg13g2_dfrbp_1 _16915_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_01859_),
    .Q_N(_00822_),
    .Q(\dp.rf.rf[24][7] ));
 sg13g2_dfrbp_1 _16916_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01860_),
    .Q_N(_00790_),
    .Q(\dp.rf.rf[24][8] ));
 sg13g2_dfrbp_1 _16917_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01861_),
    .Q_N(_00758_),
    .Q(\dp.rf.rf[24][9] ));
 sg13g2_dfrbp_1 _16918_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01862_),
    .Q_N(_00726_),
    .Q(\dp.rf.rf[24][10] ));
 sg13g2_dfrbp_1 _16919_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(_08518_),
    .D(_01863_),
    .Q_N(_00694_),
    .Q(\dp.rf.rf[24][11] ));
 sg13g2_dfrbp_1 _16920_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_08518_),
    .D(_01864_),
    .Q_N(_00662_),
    .Q(\dp.rf.rf[24][12] ));
 sg13g2_dfrbp_1 _16921_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(_08518_),
    .D(_01865_),
    .Q_N(_00630_),
    .Q(\dp.rf.rf[24][13] ));
 sg13g2_dfrbp_1 _16922_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(_08518_),
    .D(_01866_),
    .Q_N(_00598_),
    .Q(\dp.rf.rf[24][14] ));
 sg13g2_dfrbp_1 _16923_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01867_),
    .Q_N(_00566_),
    .Q(\dp.rf.rf[24][15] ));
 sg13g2_dfrbp_1 _16924_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01868_),
    .Q_N(_00534_),
    .Q(\dp.rf.rf[24][16] ));
 sg13g2_dfrbp_1 _16925_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(_08518_),
    .D(_01869_),
    .Q_N(_00502_),
    .Q(\dp.rf.rf[24][17] ));
 sg13g2_dfrbp_1 _16926_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01870_),
    .Q_N(_00471_),
    .Q(\dp.rf.rf[24][18] ));
 sg13g2_dfrbp_1 _16927_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(_08518_),
    .D(_01871_),
    .Q_N(_00439_),
    .Q(\dp.rf.rf[24][19] ));
 sg13g2_dfrbp_1 _16928_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(_08518_),
    .D(_01872_),
    .Q_N(_00408_),
    .Q(\dp.rf.rf[24][20] ));
 sg13g2_dfrbp_1 _16929_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01873_),
    .Q_N(_00376_),
    .Q(\dp.rf.rf[24][21] ));
 sg13g2_dfrbp_1 _16930_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01874_),
    .Q_N(_00344_),
    .Q(\dp.rf.rf[24][22] ));
 sg13g2_dfrbp_1 _16931_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01875_),
    .Q_N(_00312_),
    .Q(\dp.rf.rf[24][23] ));
 sg13g2_dfrbp_1 _16932_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(_08518_),
    .D(_01876_),
    .Q_N(_00280_),
    .Q(\dp.rf.rf[24][24] ));
 sg13g2_dfrbp_1 _16933_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_01877_),
    .Q_N(_00248_),
    .Q(\dp.rf.rf[24][25] ));
 sg13g2_dfrbp_1 _16934_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01878_),
    .Q_N(_00216_),
    .Q(\dp.rf.rf[24][26] ));
 sg13g2_dfrbp_1 _16935_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01879_),
    .Q_N(_00184_),
    .Q(\dp.rf.rf[24][27] ));
 sg13g2_dfrbp_1 _16936_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01880_),
    .Q_N(_00152_),
    .Q(\dp.rf.rf[24][28] ));
 sg13g2_dfrbp_1 _16937_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01881_),
    .Q_N(_00120_),
    .Q(\dp.rf.rf[24][29] ));
 sg13g2_dfrbp_1 _16938_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01882_),
    .Q_N(_00088_),
    .Q(\dp.rf.rf[24][30] ));
 sg13g2_dfrbp_1 _16939_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01883_),
    .Q_N(_00056_),
    .Q(\dp.rf.rf[24][31] ));
 sg13g2_dfrbp_1 _16940_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_08518_),
    .D(_01884_),
    .Q_N(_00023_),
    .Q(\dp.rf.rf[23][0] ));
 sg13g2_dfrbp_1 _16941_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01885_),
    .Q_N(_01013_),
    .Q(\dp.rf.rf[23][1] ));
 sg13g2_dfrbp_1 _16942_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01886_),
    .Q_N(_00981_),
    .Q(\dp.rf.rf[23][2] ));
 sg13g2_dfrbp_1 _16943_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_01887_),
    .Q_N(_00949_),
    .Q(\dp.rf.rf[23][3] ));
 sg13g2_dfrbp_1 _16944_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01888_),
    .Q_N(_00917_),
    .Q(\dp.rf.rf[23][4] ));
 sg13g2_dfrbp_1 _16945_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_08518_),
    .D(_01889_),
    .Q_N(_00885_),
    .Q(\dp.rf.rf[23][5] ));
 sg13g2_dfrbp_1 _16946_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01890_),
    .Q_N(_00853_),
    .Q(\dp.rf.rf[23][6] ));
 sg13g2_dfrbp_1 _16947_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01891_),
    .Q_N(_00821_),
    .Q(\dp.rf.rf[23][7] ));
 sg13g2_dfrbp_1 _16948_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01892_),
    .Q_N(_00789_),
    .Q(\dp.rf.rf[23][8] ));
 sg13g2_dfrbp_1 _16949_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(_08518_),
    .D(_01893_),
    .Q_N(_00757_),
    .Q(\dp.rf.rf[23][9] ));
 sg13g2_dfrbp_1 _16950_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_08518_),
    .D(_01894_),
    .Q_N(_00725_),
    .Q(\dp.rf.rf[23][10] ));
 sg13g2_dfrbp_1 _16951_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_01895_),
    .Q_N(_00693_),
    .Q(\dp.rf.rf[23][11] ));
 sg13g2_dfrbp_1 _16952_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01896_),
    .Q_N(_00661_),
    .Q(\dp.rf.rf[23][12] ));
 sg13g2_dfrbp_1 _16953_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_08518_),
    .D(_01897_),
    .Q_N(_00629_),
    .Q(\dp.rf.rf[23][13] ));
 sg13g2_dfrbp_1 _16954_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(_08518_),
    .D(_01898_),
    .Q_N(_00597_),
    .Q(\dp.rf.rf[23][14] ));
 sg13g2_dfrbp_1 _16955_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01899_),
    .Q_N(_00565_),
    .Q(\dp.rf.rf[23][15] ));
 sg13g2_dfrbp_1 _16956_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01900_),
    .Q_N(_00533_),
    .Q(\dp.rf.rf[23][16] ));
 sg13g2_dfrbp_1 _16957_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01901_),
    .Q_N(_00501_),
    .Q(\dp.rf.rf[23][17] ));
 sg13g2_dfrbp_1 _16958_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_01902_),
    .Q_N(_00470_),
    .Q(\dp.rf.rf[23][18] ));
 sg13g2_dfrbp_1 _16959_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01903_),
    .Q_N(_00438_),
    .Q(\dp.rf.rf[23][19] ));
 sg13g2_dfrbp_1 _16960_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(_08518_),
    .D(_01904_),
    .Q_N(_00407_),
    .Q(\dp.rf.rf[23][20] ));
 sg13g2_dfrbp_1 _16961_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01905_),
    .Q_N(_00375_),
    .Q(\dp.rf.rf[23][21] ));
 sg13g2_dfrbp_1 _16962_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01906_),
    .Q_N(_00343_),
    .Q(\dp.rf.rf[23][22] ));
 sg13g2_dfrbp_1 _16963_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01907_),
    .Q_N(_00311_),
    .Q(\dp.rf.rf[23][23] ));
 sg13g2_dfrbp_1 _16964_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(_08518_),
    .D(_01908_),
    .Q_N(_00279_),
    .Q(\dp.rf.rf[23][24] ));
 sg13g2_dfrbp_1 _16965_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01909_),
    .Q_N(_00247_),
    .Q(\dp.rf.rf[23][25] ));
 sg13g2_dfrbp_1 _16966_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01910_),
    .Q_N(_00215_),
    .Q(\dp.rf.rf[23][26] ));
 sg13g2_dfrbp_1 _16967_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(_08518_),
    .D(_01911_),
    .Q_N(_00183_),
    .Q(\dp.rf.rf[23][27] ));
 sg13g2_dfrbp_1 _16968_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01912_),
    .Q_N(_00151_),
    .Q(\dp.rf.rf[23][28] ));
 sg13g2_dfrbp_1 _16969_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01913_),
    .Q_N(_00119_),
    .Q(\dp.rf.rf[23][29] ));
 sg13g2_dfrbp_1 _16970_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(_08518_),
    .D(_01914_),
    .Q_N(_00087_),
    .Q(\dp.rf.rf[23][30] ));
 sg13g2_dfrbp_1 _16971_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01915_),
    .Q_N(_00055_),
    .Q(\dp.rf.rf[23][31] ));
 sg13g2_dfrbp_1 _16972_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_01916_),
    .Q_N(_00031_),
    .Q(\dp.rf.rf[31][0] ));
 sg13g2_dfrbp_1 _16973_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01917_),
    .Q_N(_01021_),
    .Q(\dp.rf.rf[31][1] ));
 sg13g2_dfrbp_1 _16974_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01918_),
    .Q_N(_00989_),
    .Q(\dp.rf.rf[31][2] ));
 sg13g2_dfrbp_1 _16975_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(_08518_),
    .D(_01919_),
    .Q_N(_00957_),
    .Q(\dp.rf.rf[31][3] ));
 sg13g2_dfrbp_1 _16976_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01920_),
    .Q_N(_00925_),
    .Q(\dp.rf.rf[31][4] ));
 sg13g2_dfrbp_1 _16977_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_08518_),
    .D(_01921_),
    .Q_N(_00893_),
    .Q(\dp.rf.rf[31][5] ));
 sg13g2_dfrbp_1 _16978_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01922_),
    .Q_N(_00861_),
    .Q(\dp.rf.rf[31][6] ));
 sg13g2_dfrbp_1 _16979_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01923_),
    .Q_N(_00829_),
    .Q(\dp.rf.rf[31][7] ));
 sg13g2_dfrbp_1 _16980_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01924_),
    .Q_N(_00797_),
    .Q(\dp.rf.rf[31][8] ));
 sg13g2_dfrbp_1 _16981_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_01925_),
    .Q_N(_00765_),
    .Q(\dp.rf.rf[31][9] ));
 sg13g2_dfrbp_1 _16982_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_08518_),
    .D(_01926_),
    .Q_N(_00733_),
    .Q(\dp.rf.rf[31][10] ));
 sg13g2_dfrbp_1 _16983_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01927_),
    .Q_N(_00701_),
    .Q(\dp.rf.rf[31][11] ));
 sg13g2_dfrbp_1 _16984_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(_08518_),
    .D(_01928_),
    .Q_N(_00669_),
    .Q(\dp.rf.rf[31][12] ));
 sg13g2_dfrbp_1 _16985_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(_08518_),
    .D(_01929_),
    .Q_N(_00637_),
    .Q(\dp.rf.rf[31][13] ));
 sg13g2_dfrbp_1 _16986_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01930_),
    .Q_N(_00605_),
    .Q(\dp.rf.rf[31][14] ));
 sg13g2_dfrbp_1 _16987_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_08518_),
    .D(_01931_),
    .Q_N(_00573_),
    .Q(\dp.rf.rf[31][15] ));
 sg13g2_dfrbp_1 _16988_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01932_),
    .Q_N(_00541_),
    .Q(\dp.rf.rf[31][16] ));
 sg13g2_dfrbp_1 _16989_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(_08518_),
    .D(_01933_),
    .Q_N(_00509_),
    .Q(\dp.rf.rf[31][17] ));
 sg13g2_dfrbp_1 _16990_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01934_),
    .Q_N(_00478_),
    .Q(\dp.rf.rf[31][18] ));
 sg13g2_dfrbp_1 _16991_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_08518_),
    .D(_01935_),
    .Q_N(_00446_),
    .Q(\dp.rf.rf[31][19] ));
 sg13g2_dfrbp_1 _16992_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(_08518_),
    .D(_01936_),
    .Q_N(_00415_),
    .Q(\dp.rf.rf[31][20] ));
 sg13g2_dfrbp_1 _16993_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01937_),
    .Q_N(_00383_),
    .Q(\dp.rf.rf[31][21] ));
 sg13g2_dfrbp_1 _16994_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01938_),
    .Q_N(_00351_),
    .Q(\dp.rf.rf[31][22] ));
 sg13g2_dfrbp_1 _16995_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01939_),
    .Q_N(_00319_),
    .Q(\dp.rf.rf[31][23] ));
 sg13g2_dfrbp_1 _16996_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(_08518_),
    .D(_01940_),
    .Q_N(_00287_),
    .Q(\dp.rf.rf[31][24] ));
 sg13g2_dfrbp_1 _16997_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01941_),
    .Q_N(_00255_),
    .Q(\dp.rf.rf[31][25] ));
 sg13g2_dfrbp_1 _16998_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(_08518_),
    .D(_01942_),
    .Q_N(_00223_),
    .Q(\dp.rf.rf[31][26] ));
 sg13g2_dfrbp_1 _16999_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(_08518_),
    .D(_01943_),
    .Q_N(_00191_),
    .Q(\dp.rf.rf[31][27] ));
 sg13g2_dfrbp_1 _17000_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_01944_),
    .Q_N(_00159_),
    .Q(\dp.rf.rf[31][28] ));
 sg13g2_dfrbp_1 _17001_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01945_),
    .Q_N(_00127_),
    .Q(\dp.rf.rf[31][29] ));
 sg13g2_dfrbp_1 _17002_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(_08518_),
    .D(_01946_),
    .Q_N(_00095_),
    .Q(\dp.rf.rf[31][30] ));
 sg13g2_dfrbp_1 _17003_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01947_),
    .Q_N(_00063_),
    .Q(\dp.rf.rf[31][31] ));
 sg13g2_dfrbp_1 _17004_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_08518_),
    .D(_01948_),
    .Q_N(_00021_),
    .Q(\dp.rf.rf[21][0] ));
 sg13g2_dfrbp_1 _17005_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(_08518_),
    .D(_01949_),
    .Q_N(_01011_),
    .Q(\dp.rf.rf[21][1] ));
 sg13g2_dfrbp_1 _17006_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(_08518_),
    .D(_01950_),
    .Q_N(_00979_),
    .Q(\dp.rf.rf[21][2] ));
 sg13g2_dfrbp_1 _17007_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_01951_),
    .Q_N(_00947_),
    .Q(\dp.rf.rf[21][3] ));
 sg13g2_dfrbp_1 _17008_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01952_),
    .Q_N(_00915_),
    .Q(\dp.rf.rf[21][4] ));
 sg13g2_dfrbp_1 _17009_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_08518_),
    .D(_01953_),
    .Q_N(_00883_),
    .Q(\dp.rf.rf[21][5] ));
 sg13g2_dfrbp_1 _17010_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(_08518_),
    .D(_01954_),
    .Q_N(_00851_),
    .Q(\dp.rf.rf[21][6] ));
 sg13g2_dfrbp_1 _17011_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01955_),
    .Q_N(_00819_),
    .Q(\dp.rf.rf[21][7] ));
 sg13g2_dfrbp_1 _17012_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_01956_),
    .Q_N(_00787_),
    .Q(\dp.rf.rf[21][8] ));
 sg13g2_dfrbp_1 _17013_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(_08518_),
    .D(_01957_),
    .Q_N(_00755_),
    .Q(\dp.rf.rf[21][9] ));
 sg13g2_dfrbp_1 _17014_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01958_),
    .Q_N(_00723_),
    .Q(\dp.rf.rf[21][10] ));
 sg13g2_dfrbp_1 _17015_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_01959_),
    .Q_N(_00691_),
    .Q(\dp.rf.rf[21][11] ));
 sg13g2_dfrbp_1 _17016_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01960_),
    .Q_N(_00659_),
    .Q(\dp.rf.rf[21][12] ));
 sg13g2_dfrbp_1 _17017_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(_08518_),
    .D(_01961_),
    .Q_N(_00627_),
    .Q(\dp.rf.rf[21][13] ));
 sg13g2_dfrbp_1 _17018_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01962_),
    .Q_N(_00595_),
    .Q(\dp.rf.rf[21][14] ));
 sg13g2_dfrbp_1 _17019_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(_08518_),
    .D(_01963_),
    .Q_N(_00563_),
    .Q(\dp.rf.rf[21][15] ));
 sg13g2_dfrbp_1 _17020_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(_08518_),
    .D(_01964_),
    .Q_N(_00531_),
    .Q(\dp.rf.rf[21][16] ));
 sg13g2_dfrbp_1 _17021_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(_08518_),
    .D(_01965_),
    .Q_N(_00499_),
    .Q(\dp.rf.rf[21][17] ));
 sg13g2_dfrbp_1 _17022_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01966_),
    .Q_N(_00468_),
    .Q(\dp.rf.rf[21][18] ));
 sg13g2_dfrbp_1 _17023_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_01967_),
    .Q_N(_00436_),
    .Q(\dp.rf.rf[21][19] ));
 sg13g2_dfrbp_1 _17024_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(_08518_),
    .D(_01968_),
    .Q_N(_00405_),
    .Q(\dp.rf.rf[21][20] ));
 sg13g2_dfrbp_1 _17025_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(_08518_),
    .D(_01969_),
    .Q_N(_00373_),
    .Q(\dp.rf.rf[21][21] ));
 sg13g2_dfrbp_1 _17026_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(_08518_),
    .D(_01970_),
    .Q_N(_00341_),
    .Q(\dp.rf.rf[21][22] ));
 sg13g2_dfrbp_1 _17027_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01971_),
    .Q_N(_00309_),
    .Q(\dp.rf.rf[21][23] ));
 sg13g2_dfrbp_1 _17028_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(_08518_),
    .D(_01972_),
    .Q_N(_00277_),
    .Q(\dp.rf.rf[21][24] ));
 sg13g2_dfrbp_1 _17029_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01973_),
    .Q_N(_00245_),
    .Q(\dp.rf.rf[21][25] ));
 sg13g2_dfrbp_1 _17030_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(_08518_),
    .D(_01974_),
    .Q_N(_00213_),
    .Q(\dp.rf.rf[21][26] ));
 sg13g2_dfrbp_1 _17031_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(_08518_),
    .D(_01975_),
    .Q_N(_00181_),
    .Q(\dp.rf.rf[21][27] ));
 sg13g2_dfrbp_1 _17032_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01976_),
    .Q_N(_00149_),
    .Q(\dp.rf.rf[21][28] ));
 sg13g2_dfrbp_1 _17033_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(_08518_),
    .D(_01977_),
    .Q_N(_00117_),
    .Q(\dp.rf.rf[21][29] ));
 sg13g2_dfrbp_1 _17034_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_01978_),
    .Q_N(_00085_),
    .Q(\dp.rf.rf[21][30] ));
 sg13g2_dfrbp_1 _17035_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_01979_),
    .Q_N(_00053_),
    .Q(\dp.rf.rf[21][31] ));
 sg13g2_dfrbp_1 _17036_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(_08518_),
    .D(_01980_),
    .Q_N(_00006_),
    .Q(\dp.rf.rf[6][0] ));
 sg13g2_dfrbp_1 _17037_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_08518_),
    .D(_01981_),
    .Q_N(_00996_),
    .Q(\dp.rf.rf[6][1] ));
 sg13g2_dfrbp_1 _17038_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(_08518_),
    .D(_01982_),
    .Q_N(_00964_),
    .Q(\dp.rf.rf[6][2] ));
 sg13g2_dfrbp_1 _17039_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(_08518_),
    .D(_01983_),
    .Q_N(_00932_),
    .Q(\dp.rf.rf[6][3] ));
 sg13g2_dfrbp_1 _17040_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(_01984_),
    .Q_N(_00900_),
    .Q(\dp.rf.rf[6][4] ));
 sg13g2_dfrbp_1 _17041_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_08518_),
    .D(_01985_),
    .Q_N(_00868_),
    .Q(\dp.rf.rf[6][5] ));
 sg13g2_dfrbp_1 _17042_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_08518_),
    .D(_01986_),
    .Q_N(_00836_),
    .Q(\dp.rf.rf[6][6] ));
 sg13g2_dfrbp_1 _17043_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_01987_),
    .Q_N(_00804_),
    .Q(\dp.rf.rf[6][7] ));
 sg13g2_dfrbp_1 _17044_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_01988_),
    .Q_N(_00772_),
    .Q(\dp.rf.rf[6][8] ));
 sg13g2_dfrbp_1 _17045_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_01989_),
    .Q_N(_00740_),
    .Q(\dp.rf.rf[6][9] ));
 sg13g2_dfrbp_1 _17046_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(_08518_),
    .D(_01990_),
    .Q_N(_00708_),
    .Q(\dp.rf.rf[6][10] ));
 sg13g2_dfrbp_1 _17047_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_01991_),
    .Q_N(_00676_),
    .Q(\dp.rf.rf[6][11] ));
 sg13g2_dfrbp_1 _17048_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_01992_),
    .Q_N(_00644_),
    .Q(\dp.rf.rf[6][12] ));
 sg13g2_dfrbp_1 _17049_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_01993_),
    .Q_N(_00612_),
    .Q(\dp.rf.rf[6][13] ));
 sg13g2_dfrbp_1 _17050_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_01994_),
    .Q_N(_00580_),
    .Q(\dp.rf.rf[6][14] ));
 sg13g2_dfrbp_1 _17051_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_01995_),
    .Q_N(_00548_),
    .Q(\dp.rf.rf[6][15] ));
 sg13g2_dfrbp_1 _17052_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_01996_),
    .Q_N(_00516_),
    .Q(\dp.rf.rf[6][16] ));
 sg13g2_dfrbp_1 _17053_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(_08518_),
    .D(_01997_),
    .Q_N(_00484_),
    .Q(\dp.rf.rf[6][17] ));
 sg13g2_dfrbp_1 _17054_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(_08518_),
    .D(_01998_),
    .Q_N(_00453_),
    .Q(\dp.rf.rf[6][18] ));
 sg13g2_dfrbp_1 _17055_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_01999_),
    .Q_N(_00421_),
    .Q(\dp.rf.rf[6][19] ));
 sg13g2_dfrbp_1 _17056_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_02000_),
    .Q_N(_00390_),
    .Q(\dp.rf.rf[6][20] ));
 sg13g2_dfrbp_1 _17057_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_02001_),
    .Q_N(_00358_),
    .Q(\dp.rf.rf[6][21] ));
 sg13g2_dfrbp_1 _17058_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(_08518_),
    .D(_02002_),
    .Q_N(_00326_),
    .Q(\dp.rf.rf[6][22] ));
 sg13g2_dfrbp_1 _17059_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(_08518_),
    .D(_02003_),
    .Q_N(_00294_),
    .Q(\dp.rf.rf[6][23] ));
 sg13g2_dfrbp_1 _17060_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_02004_),
    .Q_N(_00262_),
    .Q(\dp.rf.rf[6][24] ));
 sg13g2_dfrbp_1 _17061_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_02005_),
    .Q_N(_00230_),
    .Q(\dp.rf.rf[6][25] ));
 sg13g2_dfrbp_1 _17062_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_02006_),
    .Q_N(_00198_),
    .Q(\dp.rf.rf[6][26] ));
 sg13g2_dfrbp_1 _17063_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_02007_),
    .Q_N(_00166_),
    .Q(\dp.rf.rf[6][27] ));
 sg13g2_dfrbp_1 _17064_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_02008_),
    .Q_N(_00134_),
    .Q(\dp.rf.rf[6][28] ));
 sg13g2_dfrbp_1 _17065_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_02009_),
    .Q_N(_00102_),
    .Q(\dp.rf.rf[6][29] ));
 sg13g2_dfrbp_1 _17066_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_02010_),
    .Q_N(_00070_),
    .Q(\dp.rf.rf[6][30] ));
 sg13g2_dfrbp_1 _17067_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_02011_),
    .Q_N(_00038_),
    .Q(\dp.rf.rf[6][31] ));
 sg13g2_dfrbp_1 _17068_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_08518_),
    .D(_02012_),
    .Q_N(_00005_),
    .Q(\dp.rf.rf[5][0] ));
 sg13g2_dfrbp_1 _17069_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_08518_),
    .D(_02013_),
    .Q_N(_00995_),
    .Q(\dp.rf.rf[5][1] ));
 sg13g2_dfrbp_1 _17070_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_02014_),
    .Q_N(_00963_),
    .Q(\dp.rf.rf[5][2] ));
 sg13g2_dfrbp_1 _17071_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(_08518_),
    .D(_02015_),
    .Q_N(_00931_),
    .Q(\dp.rf.rf[5][3] ));
 sg13g2_dfrbp_1 _17072_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(_08518_),
    .D(_02016_),
    .Q_N(_00899_),
    .Q(\dp.rf.rf[5][4] ));
 sg13g2_dfrbp_1 _17073_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(_08518_),
    .D(_02017_),
    .Q_N(_00867_),
    .Q(\dp.rf.rf[5][5] ));
 sg13g2_dfrbp_1 _17074_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_08518_),
    .D(_02018_),
    .Q_N(_00835_),
    .Q(\dp.rf.rf[5][6] ));
 sg13g2_dfrbp_1 _17075_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_02019_),
    .Q_N(_00803_),
    .Q(\dp.rf.rf[5][7] ));
 sg13g2_dfrbp_1 _17076_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_02020_),
    .Q_N(_00771_),
    .Q(\dp.rf.rf[5][8] ));
 sg13g2_dfrbp_1 _17077_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(_08518_),
    .D(_02021_),
    .Q_N(_00739_),
    .Q(\dp.rf.rf[5][9] ));
 sg13g2_dfrbp_1 _17078_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(_08518_),
    .D(_02022_),
    .Q_N(_00707_),
    .Q(\dp.rf.rf[5][10] ));
 sg13g2_dfrbp_1 _17079_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(_08518_),
    .D(_02023_),
    .Q_N(_00675_),
    .Q(\dp.rf.rf[5][11] ));
 sg13g2_dfrbp_1 _17080_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(_08518_),
    .D(_02024_),
    .Q_N(_00643_),
    .Q(\dp.rf.rf[5][12] ));
 sg13g2_dfrbp_1 _17081_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(_08518_),
    .D(_02025_),
    .Q_N(_00611_),
    .Q(\dp.rf.rf[5][13] ));
 sg13g2_dfrbp_1 _17082_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_02026_),
    .Q_N(_00579_),
    .Q(\dp.rf.rf[5][14] ));
 sg13g2_dfrbp_1 _17083_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(_08518_),
    .D(_02027_),
    .Q_N(_00547_),
    .Q(\dp.rf.rf[5][15] ));
 sg13g2_dfrbp_1 _17084_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_02028_),
    .Q_N(_00515_),
    .Q(\dp.rf.rf[5][16] ));
 sg13g2_dfrbp_1 _17085_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(_08518_),
    .D(_02029_),
    .Q_N(_00483_),
    .Q(\dp.rf.rf[5][17] ));
 sg13g2_dfrbp_1 _17086_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(_08518_),
    .D(_02030_),
    .Q_N(_00452_),
    .Q(\dp.rf.rf[5][18] ));
 sg13g2_dfrbp_1 _17087_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_02031_),
    .Q_N(_00420_),
    .Q(\dp.rf.rf[5][19] ));
 sg13g2_dfrbp_1 _17088_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(_08518_),
    .D(_02032_),
    .Q_N(_00389_),
    .Q(\dp.rf.rf[5][20] ));
 sg13g2_dfrbp_1 _17089_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_02033_),
    .Q_N(_00357_),
    .Q(\dp.rf.rf[5][21] ));
 sg13g2_dfrbp_1 _17090_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(_08518_),
    .D(_02034_),
    .Q_N(_00325_),
    .Q(\dp.rf.rf[5][22] ));
 sg13g2_dfrbp_1 _17091_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(_08518_),
    .D(_02035_),
    .Q_N(_00293_),
    .Q(\dp.rf.rf[5][23] ));
 sg13g2_dfrbp_1 _17092_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(_08518_),
    .D(_02036_),
    .Q_N(_00261_),
    .Q(\dp.rf.rf[5][24] ));
 sg13g2_dfrbp_1 _17093_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_02037_),
    .Q_N(_00229_),
    .Q(\dp.rf.rf[5][25] ));
 sg13g2_dfrbp_1 _17094_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(_08518_),
    .D(_02038_),
    .Q_N(_00197_),
    .Q(\dp.rf.rf[5][26] ));
 sg13g2_dfrbp_1 _17095_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_02039_),
    .Q_N(_00165_),
    .Q(\dp.rf.rf[5][27] ));
 sg13g2_dfrbp_1 _17096_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(_08518_),
    .D(_02040_),
    .Q_N(_00133_),
    .Q(\dp.rf.rf[5][28] ));
 sg13g2_dfrbp_1 _17097_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_02041_),
    .Q_N(_00101_),
    .Q(\dp.rf.rf[5][29] ));
 sg13g2_dfrbp_1 _17098_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_02042_),
    .Q_N(_00069_),
    .Q(\dp.rf.rf[5][30] ));
 sg13g2_dfrbp_1 _17099_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(_08518_),
    .D(_02043_),
    .Q_N(_00037_),
    .Q(\dp.rf.rf[5][31] ));
 sg13g2_dfrbp_1 _17100_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net955),
    .D(_02044_),
    .Q_N(_01022_),
    .Q(net100));
 sg13g2_dfrbp_1 _17101_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net955),
    .D(_02045_),
    .Q_N(_01023_),
    .Q(net111));
 sg13g2_dfrbp_1 _17102_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(_08518_),
    .D(_02046_),
    .Q_N(_00003_),
    .Q(\dp.rf.rf[3][0] ));
 sg13g2_dfrbp_1 _17103_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_02047_),
    .Q_N(_00993_),
    .Q(\dp.rf.rf[3][1] ));
 sg13g2_dfrbp_1 _17104_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_02048_),
    .Q_N(_00961_),
    .Q(\dp.rf.rf[3][2] ));
 sg13g2_dfrbp_1 _17105_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(_08518_),
    .D(_02049_),
    .Q_N(_00929_),
    .Q(\dp.rf.rf[3][3] ));
 sg13g2_dfrbp_1 _17106_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_02050_),
    .Q_N(_00897_),
    .Q(\dp.rf.rf[3][4] ));
 sg13g2_dfrbp_1 _17107_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(_08518_),
    .D(_02051_),
    .Q_N(_00865_),
    .Q(\dp.rf.rf[3][5] ));
 sg13g2_dfrbp_1 _17108_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(_08518_),
    .D(_02052_),
    .Q_N(_00833_),
    .Q(\dp.rf.rf[3][6] ));
 sg13g2_dfrbp_1 _17109_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(_08518_),
    .D(_02053_),
    .Q_N(_00801_),
    .Q(\dp.rf.rf[3][7] ));
 sg13g2_dfrbp_1 _17110_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(_08518_),
    .D(_02054_),
    .Q_N(_00769_),
    .Q(\dp.rf.rf[3][8] ));
 sg13g2_dfrbp_1 _17111_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_02055_),
    .Q_N(_00737_),
    .Q(\dp.rf.rf[3][9] ));
 sg13g2_dfrbp_1 _17112_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(_08518_),
    .D(_02056_),
    .Q_N(_00705_),
    .Q(\dp.rf.rf[3][10] ));
 sg13g2_dfrbp_1 _17113_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(_08518_),
    .D(_02057_),
    .Q_N(_00673_),
    .Q(\dp.rf.rf[3][11] ));
 sg13g2_dfrbp_1 _17114_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(_08518_),
    .D(_02058_),
    .Q_N(_00641_),
    .Q(\dp.rf.rf[3][12] ));
 sg13g2_dfrbp_1 _17115_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(_08518_),
    .D(_02059_),
    .Q_N(_00609_),
    .Q(\dp.rf.rf[3][13] ));
 sg13g2_dfrbp_1 _17116_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(_08518_),
    .D(_02060_),
    .Q_N(_00577_),
    .Q(\dp.rf.rf[3][14] ));
 sg13g2_dfrbp_1 _17117_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(_08518_),
    .D(_02061_),
    .Q_N(_00545_),
    .Q(\dp.rf.rf[3][15] ));
 sg13g2_dfrbp_1 _17118_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_02062_),
    .Q_N(_00513_),
    .Q(\dp.rf.rf[3][16] ));
 sg13g2_dfrbp_1 _17119_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(_08518_),
    .D(_02063_),
    .Q_N(_00481_),
    .Q(\dp.rf.rf[3][17] ));
 sg13g2_dfrbp_1 _17120_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(_08518_),
    .D(_02064_),
    .Q_N(_00450_),
    .Q(\dp.rf.rf[3][18] ));
 sg13g2_dfrbp_1 _17121_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_08518_),
    .D(_02065_),
    .Q_N(_00418_),
    .Q(\dp.rf.rf[3][19] ));
 sg13g2_dfrbp_1 _17122_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(_08518_),
    .D(_02066_),
    .Q_N(_00387_),
    .Q(\dp.rf.rf[3][20] ));
 sg13g2_dfrbp_1 _17123_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(_08518_),
    .D(_02067_),
    .Q_N(_00355_),
    .Q(\dp.rf.rf[3][21] ));
 sg13g2_dfrbp_1 _17124_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(_08518_),
    .D(_02068_),
    .Q_N(_00323_),
    .Q(\dp.rf.rf[3][22] ));
 sg13g2_dfrbp_1 _17125_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(_08518_),
    .D(_02069_),
    .Q_N(_00291_),
    .Q(\dp.rf.rf[3][23] ));
 sg13g2_dfrbp_1 _17126_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(_08518_),
    .D(_02070_),
    .Q_N(_00259_),
    .Q(\dp.rf.rf[3][24] ));
 sg13g2_dfrbp_1 _17127_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(_08518_),
    .D(_02071_),
    .Q_N(_00227_),
    .Q(\dp.rf.rf[3][25] ));
 sg13g2_dfrbp_1 _17128_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(_08518_),
    .D(_02072_),
    .Q_N(_00195_),
    .Q(\dp.rf.rf[3][26] ));
 sg13g2_dfrbp_1 _17129_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(_08518_),
    .D(_02073_),
    .Q_N(_00163_),
    .Q(\dp.rf.rf[3][27] ));
 sg13g2_dfrbp_1 _17130_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(_08518_),
    .D(_02074_),
    .Q_N(_00131_),
    .Q(\dp.rf.rf[3][28] ));
 sg13g2_dfrbp_1 _17131_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(_08518_),
    .D(_02075_),
    .Q_N(_00099_),
    .Q(\dp.rf.rf[3][29] ));
 sg13g2_dfrbp_1 _17132_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(_08518_),
    .D(_02076_),
    .Q_N(_00067_),
    .Q(\dp.rf.rf[3][30] ));
 sg13g2_dfrbp_1 _17133_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(_08518_),
    .D(_02077_),
    .Q_N(_00035_),
    .Q(\dp.rf.rf[3][31] ));
 sg13g2_tiehi _17134_ ();
 sg13g2_buf_2 fanout1164 (.A(net1166),
    .X(net1164));
 sg13g2_buf_2 fanout1165 (.A(net1166),
    .X(net1165));
 sg13g2_buf_1 fanout1166 (.A(net1177),
    .X(net1166));
 sg13g2_buf_2 fanout1167 (.A(net1168),
    .X(net1167));
 sg13g2_buf_4 fanout1168 (.X(net1168),
    .A(net1169));
 sg13g2_buf_4 fanout1169 (.X(net1169),
    .A(net1177));
 sg13g2_buf_2 fanout1170 (.A(net1174),
    .X(net1170));
 sg13g2_buf_1 fanout1171 (.A(net1174),
    .X(net1171));
 sg13g2_buf_2 fanout1172 (.A(net1174),
    .X(net1172));
 sg13g2_buf_1 fanout1173 (.A(net1174),
    .X(net1173));
 sg13g2_buf_1 fanout1174 (.A(net1177),
    .X(net1174));
 sg13g2_buf_2 fanout1175 (.A(net1177),
    .X(net1175));
 sg13g2_buf_2 fanout1176 (.A(net1177),
    .X(net1176));
 sg13g2_buf_2 fanout1177 (.A(net1203),
    .X(net1177));
 sg13g2_buf_4 fanout1178 (.X(net1178),
    .A(net1180));
 sg13g2_buf_4 fanout1179 (.X(net1179),
    .A(net1181));
 sg13g2_buf_1 fanout1180 (.A(net1181),
    .X(net1180));
 sg13g2_buf_4 fanout1181 (.X(net1181),
    .A(net1203));
 sg13g2_buf_4 fanout1182 (.X(net1182),
    .A(net1184));
 sg13g2_buf_1 fanout1183 (.A(net1184),
    .X(net1183));
 sg13g2_buf_2 fanout1184 (.A(net1187),
    .X(net1184));
 sg13g2_buf_2 fanout1185 (.A(net1186),
    .X(net1185));
 sg13g2_buf_4 fanout1186 (.X(net1186),
    .A(net1187));
 sg13g2_buf_2 fanout1187 (.A(net1203),
    .X(net1187));
 sg13g2_buf_4 fanout1188 (.X(net1188),
    .A(net1189));
 sg13g2_buf_2 fanout1189 (.A(net1190),
    .X(net1189));
 sg13g2_buf_1 fanout1190 (.A(net1203),
    .X(net1190));
 sg13g2_buf_2 fanout1191 (.A(net1193),
    .X(net1191));
 sg13g2_buf_1 fanout1192 (.A(net1193),
    .X(net1192));
 sg13g2_buf_2 fanout1193 (.A(net1202),
    .X(net1193));
 sg13g2_buf_2 fanout1194 (.A(net1197),
    .X(net1194));
 sg13g2_buf_2 fanout1195 (.A(net1197),
    .X(net1195));
 sg13g2_buf_4 fanout1196 (.X(net1196),
    .A(net1197));
 sg13g2_buf_1 fanout1197 (.A(net1202),
    .X(net1197));
 sg13g2_buf_2 fanout1198 (.A(net1199),
    .X(net1198));
 sg13g2_buf_2 fanout1199 (.A(net1202),
    .X(net1199));
 sg13g2_buf_4 fanout1200 (.X(net1200),
    .A(net1202));
 sg13g2_buf_2 fanout1201 (.A(net1202),
    .X(net1201));
 sg13g2_buf_2 fanout1202 (.A(net1203),
    .X(net1202));
 sg13g2_buf_2 fanout1203 (.A(net1204),
    .X(net1203));
 sg13g2_buf_1 fanout1204 (.A(net8),
    .X(net1204));
 sg13g2_buf_4 fanout1205 (.X(net1205),
    .A(net1206));
 sg13g2_buf_4 fanout1206 (.X(net1206),
    .A(net1210));
 sg13g2_buf_2 fanout1207 (.A(net1209),
    .X(net1207));
 sg13g2_buf_2 fanout1208 (.A(net1209),
    .X(net1208));
 sg13g2_buf_2 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_2 fanout1210 (.A(net1224),
    .X(net1210));
 sg13g2_buf_2 fanout1211 (.A(net1215),
    .X(net1211));
 sg13g2_buf_2 fanout1212 (.A(net1215),
    .X(net1212));
 sg13g2_buf_2 fanout1213 (.A(net1215),
    .X(net1213));
 sg13g2_buf_2 fanout1214 (.A(net1215),
    .X(net1214));
 sg13g2_buf_1 fanout1215 (.A(net1224),
    .X(net1215));
 sg13g2_buf_2 fanout1216 (.A(net1218),
    .X(net1216));
 sg13g2_buf_2 fanout1217 (.A(net1218),
    .X(net1217));
 sg13g2_buf_2 fanout1218 (.A(net1224),
    .X(net1218));
 sg13g2_buf_2 fanout1219 (.A(net1220),
    .X(net1219));
 sg13g2_buf_2 fanout1220 (.A(net1221),
    .X(net1220));
 sg13g2_buf_2 fanout1221 (.A(net1224),
    .X(net1221));
 sg13g2_buf_4 fanout1222 (.X(net1222),
    .A(net1223));
 sg13g2_buf_1 fanout1223 (.A(net1224),
    .X(net1223));
 sg13g2_buf_1 fanout1224 (.A(net1236),
    .X(net1224));
 sg13g2_buf_4 fanout1225 (.X(net1225),
    .A(net1226));
 sg13g2_buf_4 fanout1226 (.X(net1226),
    .A(net1231));
 sg13g2_buf_2 fanout1227 (.A(net1228),
    .X(net1227));
 sg13g2_buf_2 fanout1228 (.A(net1231),
    .X(net1228));
 sg13g2_buf_4 fanout1229 (.X(net1229),
    .A(net1231));
 sg13g2_buf_2 fanout1230 (.A(net1231),
    .X(net1230));
 sg13g2_buf_2 fanout1231 (.A(net1236),
    .X(net1231));
 sg13g2_buf_2 fanout1232 (.A(net1233),
    .X(net1232));
 sg13g2_buf_2 fanout1233 (.A(net1236),
    .X(net1233));
 sg13g2_buf_2 fanout1234 (.A(net1235),
    .X(net1234));
 sg13g2_buf_2 fanout1235 (.A(net1236),
    .X(net1235));
 sg13g2_buf_1 fanout1236 (.A(net7),
    .X(net1236));
 sg13g2_buf_2 fanout1237 (.A(net1238),
    .X(net1237));
 sg13g2_buf_2 fanout1238 (.A(net6),
    .X(net1238));
 sg13g2_buf_2 fanout1239 (.A(net1240),
    .X(net1239));
 sg13g2_buf_1 fanout1240 (.A(net1241),
    .X(net1240));
 sg13g2_buf_1 fanout1241 (.A(net5),
    .X(net1241));
 sg13g2_buf_2 fanout1242 (.A(net4),
    .X(net1242));
 sg13g2_buf_1 fanout1243 (.A(net4),
    .X(net1243));
 sg13g2_buf_2 fanout1244 (.A(net32),
    .X(net1244));
 sg13g2_buf_2 fanout1245 (.A(net1246),
    .X(net1245));
 sg13g2_buf_1 fanout1246 (.A(net30),
    .X(net1246));
 sg13g2_buf_2 fanout1247 (.A(net3),
    .X(net1247));
 sg13g2_buf_2 fanout1248 (.A(net29),
    .X(net1248));
 sg13g2_buf_2 fanout1249 (.A(net1250),
    .X(net1249));
 sg13g2_buf_1 fanout1250 (.A(net28),
    .X(net1250));
 sg13g2_buf_2 fanout1251 (.A(net26),
    .X(net1251));
 sg13g2_buf_1 fanout1252 (.A(net26),
    .X(net1252));
 sg13g2_buf_2 fanout1253 (.A(net24),
    .X(net1253));
 sg13g2_buf_2 fanout1254 (.A(net23),
    .X(net1254));
 sg13g2_buf_1 fanout1255 (.A(net23),
    .X(net1255));
 sg13g2_buf_2 fanout1256 (.A(net1257),
    .X(net1256));
 sg13g2_buf_1 fanout1257 (.A(net2),
    .X(net1257));
 sg13g2_buf_2 fanout1258 (.A(net1261),
    .X(net1258));
 sg13g2_buf_1 fanout1259 (.A(net1261),
    .X(net1259));
 sg13g2_buf_2 fanout1260 (.A(net1261),
    .X(net1260));
 sg13g2_buf_2 fanout1261 (.A(net17),
    .X(net1261));
 sg13g2_buf_2 fanout1262 (.A(net1264),
    .X(net1262));
 sg13g2_buf_2 fanout1263 (.A(net1264),
    .X(net1263));
 sg13g2_buf_2 fanout1264 (.A(net1274),
    .X(net1264));
 sg13g2_buf_2 fanout1265 (.A(net1274),
    .X(net1265));
 sg13g2_buf_2 fanout1266 (.A(net1268),
    .X(net1266));
 sg13g2_buf_1 fanout1267 (.A(net1268),
    .X(net1267));
 sg13g2_buf_2 fanout1268 (.A(net1269),
    .X(net1268));
 sg13g2_buf_2 fanout1269 (.A(net1274),
    .X(net1269));
 sg13g2_buf_2 fanout1270 (.A(net1272),
    .X(net1270));
 sg13g2_buf_2 fanout1271 (.A(net1272),
    .X(net1271));
 sg13g2_buf_2 fanout1272 (.A(net1273),
    .X(net1272));
 sg13g2_buf_2 fanout1273 (.A(net1274),
    .X(net1273));
 sg13g2_buf_2 fanout1274 (.A(net16),
    .X(net1274));
 sg13g2_buf_2 fanout1275 (.A(net1277),
    .X(net1275));
 sg13g2_buf_2 fanout1276 (.A(net1277),
    .X(net1276));
 sg13g2_buf_2 fanout1277 (.A(net15),
    .X(net1277));
 sg13g2_buf_4 fanout1278 (.X(net1278),
    .A(net1279));
 sg13g2_buf_1 fanout1279 (.A(net1281),
    .X(net1279));
 sg13g2_buf_4 fanout1280 (.X(net1280),
    .A(net1281));
 sg13g2_buf_1 fanout1281 (.A(net1302),
    .X(net1281));
 sg13g2_buf_4 fanout1282 (.X(net1282),
    .A(net1285));
 sg13g2_buf_2 fanout1283 (.A(net1285),
    .X(net1283));
 sg13g2_buf_2 fanout1284 (.A(net1285),
    .X(net1284));
 sg13g2_buf_2 fanout1285 (.A(net1302),
    .X(net1285));
 sg13g2_buf_4 fanout1286 (.X(net1286),
    .A(net1290));
 sg13g2_buf_2 fanout1287 (.A(net1290),
    .X(net1287));
 sg13g2_buf_4 fanout1288 (.X(net1288),
    .A(net1289));
 sg13g2_buf_4 fanout1289 (.X(net1289),
    .A(net1290));
 sg13g2_buf_2 fanout1290 (.A(net1302),
    .X(net1290));
 sg13g2_buf_4 fanout1291 (.X(net1291),
    .A(net1292));
 sg13g2_buf_2 fanout1292 (.A(net1302),
    .X(net1292));
 sg13g2_buf_2 fanout1293 (.A(net1296),
    .X(net1293));
 sg13g2_buf_1 fanout1294 (.A(net1296),
    .X(net1294));
 sg13g2_buf_4 fanout1295 (.X(net1295),
    .A(net1296));
 sg13g2_buf_2 fanout1296 (.A(net1302),
    .X(net1296));
 sg13g2_buf_2 fanout1297 (.A(net1300),
    .X(net1297));
 sg13g2_buf_2 fanout1298 (.A(net1300),
    .X(net1298));
 sg13g2_buf_2 fanout1299 (.A(net1300),
    .X(net1299));
 sg13g2_buf_1 fanout1300 (.A(net1301),
    .X(net1300));
 sg13g2_buf_2 fanout1301 (.A(net1302),
    .X(net1301));
 sg13g2_buf_2 fanout1302 (.A(net14),
    .X(net1302));
 sg13g2_buf_2 fanout1303 (.A(net1305),
    .X(net1303));
 sg13g2_buf_1 fanout1304 (.A(net1305),
    .X(net1304));
 sg13g2_buf_2 fanout1305 (.A(net1314),
    .X(net1305));
 sg13g2_buf_4 fanout1306 (.X(net1306),
    .A(net1314));
 sg13g2_buf_4 fanout1307 (.X(net1307),
    .A(net1314));
 sg13g2_buf_2 fanout1308 (.A(net1310),
    .X(net1308));
 sg13g2_buf_2 fanout1309 (.A(net1310),
    .X(net1309));
 sg13g2_buf_4 fanout1310 (.X(net1310),
    .A(net1313));
 sg13g2_buf_4 fanout1311 (.X(net1311),
    .A(net1313));
 sg13g2_buf_4 fanout1312 (.X(net1312),
    .A(net1313));
 sg13g2_buf_2 fanout1313 (.A(net1314),
    .X(net1313));
 sg13g2_buf_1 fanout1314 (.A(net1345),
    .X(net1314));
 sg13g2_buf_2 fanout1315 (.A(net1318),
    .X(net1315));
 sg13g2_buf_2 fanout1316 (.A(net1317),
    .X(net1316));
 sg13g2_buf_2 fanout1317 (.A(net1318),
    .X(net1317));
 sg13g2_buf_2 fanout1318 (.A(net1329),
    .X(net1318));
 sg13g2_buf_2 fanout1319 (.A(net1323),
    .X(net1319));
 sg13g2_buf_2 fanout1320 (.A(net1323),
    .X(net1320));
 sg13g2_buf_2 fanout1321 (.A(net1323),
    .X(net1321));
 sg13g2_buf_1 fanout1322 (.A(net1323),
    .X(net1322));
 sg13g2_buf_1 fanout1323 (.A(net1329),
    .X(net1323));
 sg13g2_buf_2 fanout1324 (.A(net1325),
    .X(net1324));
 sg13g2_buf_4 fanout1325 (.X(net1325),
    .A(net1329));
 sg13g2_buf_4 fanout1326 (.X(net1326),
    .A(net1328));
 sg13g2_buf_2 fanout1327 (.A(net1328),
    .X(net1327));
 sg13g2_buf_2 fanout1328 (.A(net1329),
    .X(net1328));
 sg13g2_buf_1 fanout1329 (.A(net1345),
    .X(net1329));
 sg13g2_buf_4 fanout1330 (.X(net1330),
    .A(net1333));
 sg13g2_buf_2 fanout1331 (.A(net1332),
    .X(net1331));
 sg13g2_buf_2 fanout1332 (.A(net1333),
    .X(net1332));
 sg13g2_buf_2 fanout1333 (.A(net1339),
    .X(net1333));
 sg13g2_buf_2 fanout1334 (.A(net1335),
    .X(net1334));
 sg13g2_buf_4 fanout1335 (.X(net1335),
    .A(net1339));
 sg13g2_buf_2 fanout1336 (.A(net1337),
    .X(net1336));
 sg13g2_buf_4 fanout1337 (.X(net1337),
    .A(net1338));
 sg13g2_buf_4 fanout1338 (.X(net1338),
    .A(net1339));
 sg13g2_buf_1 fanout1339 (.A(net1345),
    .X(net1339));
 sg13g2_buf_2 fanout1340 (.A(net1341),
    .X(net1340));
 sg13g2_buf_2 fanout1341 (.A(net1344),
    .X(net1341));
 sg13g2_buf_2 fanout1342 (.A(net1343),
    .X(net1342));
 sg13g2_buf_2 fanout1343 (.A(net1344),
    .X(net1343));
 sg13g2_buf_2 fanout1344 (.A(net1345),
    .X(net1344));
 sg13g2_buf_1 fanout1345 (.A(net1390),
    .X(net1345));
 sg13g2_buf_4 fanout1346 (.X(net1346),
    .A(net1350));
 sg13g2_buf_1 fanout1347 (.A(net1350),
    .X(net1347));
 sg13g2_buf_2 fanout1348 (.A(net1350),
    .X(net1348));
 sg13g2_buf_2 fanout1349 (.A(net1350),
    .X(net1349));
 sg13g2_buf_1 fanout1350 (.A(net1370),
    .X(net1350));
 sg13g2_buf_2 fanout1351 (.A(net1354),
    .X(net1351));
 sg13g2_buf_2 fanout1352 (.A(net1354),
    .X(net1352));
 sg13g2_buf_4 fanout1353 (.X(net1353),
    .A(net1354));
 sg13g2_buf_2 fanout1354 (.A(net1370),
    .X(net1354));
 sg13g2_buf_4 fanout1355 (.X(net1355),
    .A(net1356));
 sg13g2_buf_4 fanout1356 (.X(net1356),
    .A(net1359));
 sg13g2_buf_4 fanout1357 (.X(net1357),
    .A(net1358));
 sg13g2_buf_4 fanout1358 (.X(net1358),
    .A(net1359));
 sg13g2_buf_2 fanout1359 (.A(net1370),
    .X(net1359));
 sg13g2_buf_4 fanout1360 (.X(net1360),
    .A(net1369));
 sg13g2_buf_2 fanout1361 (.A(net1369),
    .X(net1361));
 sg13g2_buf_2 fanout1362 (.A(net1363),
    .X(net1362));
 sg13g2_buf_2 fanout1363 (.A(net1369),
    .X(net1363));
 sg13g2_buf_4 fanout1364 (.X(net1364),
    .A(net1369));
 sg13g2_buf_4 fanout1365 (.X(net1365),
    .A(net1369));
 sg13g2_buf_2 fanout1366 (.A(net1367),
    .X(net1366));
 sg13g2_buf_2 fanout1367 (.A(net1368),
    .X(net1367));
 sg13g2_buf_4 fanout1368 (.X(net1368),
    .A(net1369));
 sg13g2_buf_2 fanout1369 (.A(net1370),
    .X(net1369));
 sg13g2_buf_1 fanout1370 (.A(net1390),
    .X(net1370));
 sg13g2_buf_2 fanout1371 (.A(net1375),
    .X(net1371));
 sg13g2_buf_1 fanout1372 (.A(net1375),
    .X(net1372));
 sg13g2_buf_2 fanout1373 (.A(net1374),
    .X(net1373));
 sg13g2_buf_1 fanout1374 (.A(net1375),
    .X(net1374));
 sg13g2_buf_2 fanout1375 (.A(net1390),
    .X(net1375));
 sg13g2_buf_2 fanout1376 (.A(net1377),
    .X(net1376));
 sg13g2_buf_2 fanout1377 (.A(net1389),
    .X(net1377));
 sg13g2_buf_2 fanout1378 (.A(net1379),
    .X(net1378));
 sg13g2_buf_4 fanout1379 (.X(net1379),
    .A(net1381));
 sg13g2_buf_4 fanout1380 (.X(net1380),
    .A(net1381));
 sg13g2_buf_1 fanout1381 (.A(net1389),
    .X(net1381));
 sg13g2_buf_2 fanout1382 (.A(net1383),
    .X(net1382));
 sg13g2_buf_2 fanout1383 (.A(net1387),
    .X(net1383));
 sg13g2_buf_2 fanout1384 (.A(net1387),
    .X(net1384));
 sg13g2_buf_1 fanout1385 (.A(net1387),
    .X(net1385));
 sg13g2_buf_4 fanout1386 (.X(net1386),
    .A(net1387));
 sg13g2_buf_1 fanout1387 (.A(net1389),
    .X(net1387));
 sg13g2_buf_2 fanout1388 (.A(net1389),
    .X(net1388));
 sg13g2_buf_1 fanout1389 (.A(net1390),
    .X(net1389));
 sg13g2_buf_1 fanout1390 (.A(net13),
    .X(net1390));
 sg13g2_buf_2 fanout1391 (.A(net1392),
    .X(net1391));
 sg13g2_buf_2 fanout1392 (.A(net1395),
    .X(net1392));
 sg13g2_buf_2 fanout1393 (.A(net1394),
    .X(net1393));
 sg13g2_buf_2 fanout1394 (.A(net1395),
    .X(net1394));
 sg13g2_buf_2 fanout1395 (.A(net11),
    .X(net1395));
 sg13g2_buf_2 fanout1396 (.A(net1397),
    .X(net1396));
 sg13g2_buf_2 fanout1397 (.A(net1398),
    .X(net1397));
 sg13g2_buf_4 fanout1398 (.X(net1398),
    .A(net1402));
 sg13g2_buf_4 fanout1399 (.X(net1399),
    .A(net1401));
 sg13g2_buf_1 fanout1400 (.A(net1401),
    .X(net1400));
 sg13g2_buf_2 fanout1401 (.A(net1402),
    .X(net1401));
 sg13g2_buf_2 fanout1402 (.A(net10),
    .X(net1402));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_fill_8 FILLER_0_0_0 ();
 sg13g2_fill_8 FILLER_0_0_8 ();
 sg13g2_fill_8 FILLER_0_0_16 ();
 sg13g2_fill_8 FILLER_0_0_24 ();
 sg13g2_fill_8 FILLER_0_0_32 ();
 sg13g2_fill_8 FILLER_0_0_40 ();
 sg13g2_fill_8 FILLER_0_0_48 ();
 sg13g2_fill_8 FILLER_0_0_56 ();
 sg13g2_fill_8 FILLER_0_0_64 ();
 sg13g2_fill_8 FILLER_0_0_72 ();
 sg13g2_fill_8 FILLER_0_0_80 ();
 sg13g2_fill_8 FILLER_0_0_88 ();
 sg13g2_fill_8 FILLER_0_0_96 ();
 sg13g2_fill_8 FILLER_0_0_104 ();
 sg13g2_fill_8 FILLER_0_0_112 ();
 sg13g2_fill_8 FILLER_0_0_120 ();
 sg13g2_fill_8 FILLER_0_0_128 ();
 sg13g2_fill_8 FILLER_0_0_136 ();
 sg13g2_fill_8 FILLER_0_0_144 ();
 sg13g2_fill_8 FILLER_0_0_152 ();
 sg13g2_fill_8 FILLER_0_0_160 ();
 sg13g2_fill_8 FILLER_0_0_168 ();
 sg13g2_fill_8 FILLER_0_0_176 ();
 sg13g2_fill_8 FILLER_0_0_184 ();
 sg13g2_fill_8 FILLER_0_0_192 ();
 sg13g2_fill_8 FILLER_0_0_200 ();
 sg13g2_fill_4 FILLER_0_0_208 ();
 sg13g2_fill_2 FILLER_0_0_212 ();
 sg13g2_fill_1 FILLER_0_0_214 ();
 sg13g2_fill_8 FILLER_0_0_219 ();
 sg13g2_fill_8 FILLER_0_0_227 ();
 sg13g2_fill_8 FILLER_0_0_235 ();
 sg13g2_fill_8 FILLER_0_0_243 ();
 sg13g2_fill_8 FILLER_0_0_251 ();
 sg13g2_fill_8 FILLER_0_0_259 ();
 sg13g2_fill_8 FILLER_0_0_267 ();
 sg13g2_fill_8 FILLER_0_0_275 ();
 sg13g2_fill_8 FILLER_0_0_283 ();
 sg13g2_fill_8 FILLER_0_0_291 ();
 sg13g2_fill_8 FILLER_0_0_299 ();
 sg13g2_fill_8 FILLER_0_0_307 ();
 sg13g2_fill_8 FILLER_0_0_315 ();
 sg13g2_fill_8 FILLER_0_0_323 ();
 sg13g2_fill_8 FILLER_0_0_331 ();
 sg13g2_fill_8 FILLER_0_0_339 ();
 sg13g2_fill_8 FILLER_0_0_347 ();
 sg13g2_fill_8 FILLER_0_0_355 ();
 sg13g2_fill_8 FILLER_0_0_363 ();
 sg13g2_fill_8 FILLER_0_0_371 ();
 sg13g2_fill_8 FILLER_0_0_379 ();
 sg13g2_fill_8 FILLER_0_0_387 ();
 sg13g2_fill_8 FILLER_0_0_395 ();
 sg13g2_fill_8 FILLER_0_0_403 ();
 sg13g2_fill_8 FILLER_0_0_411 ();
 sg13g2_fill_8 FILLER_0_0_419 ();
 sg13g2_fill_8 FILLER_0_0_427 ();
 sg13g2_fill_8 FILLER_0_0_435 ();
 sg13g2_fill_8 FILLER_0_0_443 ();
 sg13g2_fill_8 FILLER_0_0_451 ();
 sg13g2_fill_8 FILLER_0_0_459 ();
 sg13g2_fill_8 FILLER_0_0_467 ();
 sg13g2_fill_8 FILLER_0_0_475 ();
 sg13g2_fill_8 FILLER_0_0_483 ();
 sg13g2_fill_8 FILLER_0_0_491 ();
 sg13g2_fill_8 FILLER_0_0_499 ();
 sg13g2_fill_8 FILLER_0_0_507 ();
 sg13g2_fill_8 FILLER_0_0_515 ();
 sg13g2_fill_4 FILLER_0_0_523 ();
 sg13g2_fill_1 FILLER_0_0_527 ();
 sg13g2_fill_8 FILLER_0_0_532 ();
 sg13g2_fill_8 FILLER_0_0_540 ();
 sg13g2_fill_8 FILLER_0_0_548 ();
 sg13g2_fill_8 FILLER_0_0_556 ();
 sg13g2_fill_8 FILLER_0_0_564 ();
 sg13g2_fill_8 FILLER_0_0_572 ();
 sg13g2_fill_8 FILLER_0_0_580 ();
 sg13g2_fill_8 FILLER_0_0_588 ();
 sg13g2_fill_8 FILLER_0_0_596 ();
 sg13g2_fill_8 FILLER_0_0_604 ();
 sg13g2_fill_8 FILLER_0_0_612 ();
 sg13g2_fill_8 FILLER_0_0_620 ();
 sg13g2_fill_8 FILLER_0_0_628 ();
 sg13g2_fill_8 FILLER_0_0_636 ();
 sg13g2_fill_8 FILLER_0_0_644 ();
 sg13g2_fill_8 FILLER_0_0_652 ();
 sg13g2_fill_8 FILLER_0_0_660 ();
 sg13g2_fill_8 FILLER_0_0_668 ();
 sg13g2_fill_8 FILLER_0_0_676 ();
 sg13g2_fill_8 FILLER_0_0_684 ();
 sg13g2_fill_8 FILLER_0_0_692 ();
 sg13g2_fill_1 FILLER_0_0_700 ();
 sg13g2_fill_4 FILLER_0_0_706 ();
 sg13g2_fill_2 FILLER_0_0_710 ();
 sg13g2_fill_1 FILLER_0_0_712 ();
 sg13g2_fill_8 FILLER_0_0_717 ();
 sg13g2_fill_8 FILLER_0_0_725 ();
 sg13g2_fill_8 FILLER_0_0_733 ();
 sg13g2_fill_8 FILLER_0_0_741 ();
 sg13g2_fill_8 FILLER_0_0_749 ();
 sg13g2_fill_8 FILLER_0_0_757 ();
 sg13g2_fill_8 FILLER_0_0_765 ();
 sg13g2_fill_8 FILLER_0_0_773 ();
 sg13g2_fill_8 FILLER_0_0_781 ();
 sg13g2_fill_8 FILLER_0_0_789 ();
 sg13g2_fill_8 FILLER_0_0_797 ();
 sg13g2_fill_8 FILLER_0_0_805 ();
 sg13g2_fill_8 FILLER_0_0_813 ();
 sg13g2_fill_8 FILLER_0_0_821 ();
 sg13g2_fill_8 FILLER_0_0_829 ();
 sg13g2_fill_8 FILLER_0_0_837 ();
 sg13g2_fill_8 FILLER_0_0_845 ();
 sg13g2_fill_8 FILLER_0_0_853 ();
 sg13g2_fill_8 FILLER_0_0_861 ();
 sg13g2_fill_8 FILLER_0_0_869 ();
 sg13g2_fill_8 FILLER_0_0_877 ();
 sg13g2_fill_8 FILLER_0_0_885 ();
 sg13g2_fill_8 FILLER_0_0_893 ();
 sg13g2_fill_8 FILLER_0_0_901 ();
 sg13g2_fill_8 FILLER_0_0_909 ();
 sg13g2_fill_8 FILLER_0_0_917 ();
 sg13g2_fill_8 FILLER_0_0_925 ();
 sg13g2_fill_8 FILLER_0_0_933 ();
 sg13g2_fill_8 FILLER_0_0_941 ();
 sg13g2_fill_8 FILLER_0_0_949 ();
 sg13g2_fill_8 FILLER_0_0_957 ();
 sg13g2_fill_1 FILLER_0_0_965 ();
 sg13g2_fill_8 FILLER_0_0_970 ();
 sg13g2_fill_8 FILLER_0_0_978 ();
 sg13g2_fill_8 FILLER_0_0_986 ();
 sg13g2_fill_8 FILLER_0_0_994 ();
 sg13g2_fill_2 FILLER_0_0_1002 ();
 sg13g2_fill_4 FILLER_0_0_1008 ();
 sg13g2_fill_8 FILLER_0_0_1016 ();
 sg13g2_fill_8 FILLER_0_0_1024 ();
 sg13g2_fill_8 FILLER_0_0_1032 ();
 sg13g2_fill_8 FILLER_0_0_1040 ();
 sg13g2_fill_1 FILLER_0_0_1048 ();
 sg13g2_fill_2 FILLER_0_0_1053 ();
 sg13g2_fill_2 FILLER_0_0_1059 ();
 sg13g2_fill_8 FILLER_0_0_1065 ();
 sg13g2_fill_8 FILLER_0_0_1073 ();
 sg13g2_fill_8 FILLER_0_0_1081 ();
 sg13g2_fill_8 FILLER_0_0_1089 ();
 sg13g2_fill_8 FILLER_0_0_1097 ();
 sg13g2_fill_8 FILLER_0_0_1105 ();
 sg13g2_fill_8 FILLER_0_0_1113 ();
 sg13g2_fill_8 FILLER_0_0_1121 ();
 sg13g2_fill_8 FILLER_0_0_1129 ();
 sg13g2_fill_8 FILLER_0_0_1137 ();
 sg13g2_fill_8 FILLER_0_0_1145 ();
 sg13g2_fill_8 FILLER_0_0_1153 ();
 sg13g2_fill_8 FILLER_0_0_1161 ();
 sg13g2_fill_8 FILLER_0_0_1169 ();
 sg13g2_fill_8 FILLER_0_0_1177 ();
 sg13g2_fill_8 FILLER_0_0_1185 ();
 sg13g2_fill_8 FILLER_0_0_1193 ();
 sg13g2_fill_8 FILLER_0_0_1201 ();
 sg13g2_fill_8 FILLER_0_0_1209 ();
 sg13g2_fill_8 FILLER_0_0_1217 ();
 sg13g2_fill_8 FILLER_0_0_1225 ();
 sg13g2_fill_8 FILLER_0_0_1233 ();
 sg13g2_fill_8 FILLER_0_0_1241 ();
 sg13g2_fill_8 FILLER_0_0_1249 ();
 sg13g2_fill_8 FILLER_0_0_1257 ();
 sg13g2_fill_8 FILLER_0_0_1265 ();
 sg13g2_fill_8 FILLER_0_0_1273 ();
 sg13g2_fill_8 FILLER_0_0_1281 ();
 sg13g2_fill_8 FILLER_0_0_1289 ();
 sg13g2_fill_8 FILLER_0_1_0 ();
 sg13g2_fill_8 FILLER_0_1_8 ();
 sg13g2_fill_8 FILLER_0_1_16 ();
 sg13g2_fill_8 FILLER_0_1_24 ();
 sg13g2_fill_8 FILLER_0_1_32 ();
 sg13g2_fill_8 FILLER_0_1_40 ();
 sg13g2_fill_8 FILLER_0_1_48 ();
 sg13g2_fill_8 FILLER_0_1_56 ();
 sg13g2_fill_8 FILLER_0_1_64 ();
 sg13g2_fill_8 FILLER_0_1_72 ();
 sg13g2_fill_8 FILLER_0_1_80 ();
 sg13g2_fill_8 FILLER_0_1_88 ();
 sg13g2_fill_8 FILLER_0_1_96 ();
 sg13g2_fill_8 FILLER_0_1_104 ();
 sg13g2_fill_8 FILLER_0_1_112 ();
 sg13g2_fill_8 FILLER_0_1_120 ();
 sg13g2_fill_8 FILLER_0_1_128 ();
 sg13g2_fill_8 FILLER_0_1_136 ();
 sg13g2_fill_8 FILLER_0_1_144 ();
 sg13g2_fill_8 FILLER_0_1_152 ();
 sg13g2_fill_8 FILLER_0_1_160 ();
 sg13g2_fill_8 FILLER_0_1_168 ();
 sg13g2_fill_8 FILLER_0_1_176 ();
 sg13g2_fill_8 FILLER_0_1_184 ();
 sg13g2_fill_8 FILLER_0_1_192 ();
 sg13g2_fill_8 FILLER_0_1_200 ();
 sg13g2_fill_8 FILLER_0_1_208 ();
 sg13g2_fill_8 FILLER_0_1_216 ();
 sg13g2_fill_8 FILLER_0_1_224 ();
 sg13g2_fill_8 FILLER_0_1_232 ();
 sg13g2_fill_8 FILLER_0_1_240 ();
 sg13g2_fill_8 FILLER_0_1_248 ();
 sg13g2_fill_8 FILLER_0_1_256 ();
 sg13g2_fill_8 FILLER_0_1_264 ();
 sg13g2_fill_8 FILLER_0_1_272 ();
 sg13g2_fill_8 FILLER_0_1_280 ();
 sg13g2_fill_8 FILLER_0_1_288 ();
 sg13g2_fill_8 FILLER_0_1_296 ();
 sg13g2_fill_8 FILLER_0_1_304 ();
 sg13g2_fill_8 FILLER_0_1_312 ();
 sg13g2_fill_8 FILLER_0_1_320 ();
 sg13g2_fill_8 FILLER_0_1_328 ();
 sg13g2_fill_8 FILLER_0_1_336 ();
 sg13g2_fill_8 FILLER_0_1_344 ();
 sg13g2_fill_8 FILLER_0_1_352 ();
 sg13g2_fill_8 FILLER_0_1_360 ();
 sg13g2_fill_8 FILLER_0_1_368 ();
 sg13g2_fill_8 FILLER_0_1_376 ();
 sg13g2_fill_8 FILLER_0_1_384 ();
 sg13g2_fill_8 FILLER_0_1_392 ();
 sg13g2_fill_8 FILLER_0_1_400 ();
 sg13g2_fill_8 FILLER_0_1_408 ();
 sg13g2_fill_8 FILLER_0_1_416 ();
 sg13g2_fill_8 FILLER_0_1_424 ();
 sg13g2_fill_8 FILLER_0_1_432 ();
 sg13g2_fill_8 FILLER_0_1_440 ();
 sg13g2_fill_8 FILLER_0_1_448 ();
 sg13g2_fill_8 FILLER_0_1_456 ();
 sg13g2_fill_8 FILLER_0_1_464 ();
 sg13g2_fill_8 FILLER_0_1_472 ();
 sg13g2_fill_8 FILLER_0_1_480 ();
 sg13g2_fill_8 FILLER_0_1_488 ();
 sg13g2_fill_8 FILLER_0_1_496 ();
 sg13g2_fill_8 FILLER_0_1_504 ();
 sg13g2_fill_8 FILLER_0_1_512 ();
 sg13g2_fill_8 FILLER_0_1_520 ();
 sg13g2_fill_8 FILLER_0_1_528 ();
 sg13g2_fill_4 FILLER_0_1_536 ();
 sg13g2_fill_2 FILLER_0_1_540 ();
 sg13g2_fill_2 FILLER_0_1_546 ();
 sg13g2_fill_8 FILLER_0_1_574 ();
 sg13g2_fill_4 FILLER_0_1_582 ();
 sg13g2_fill_1 FILLER_0_1_586 ();
 sg13g2_fill_8 FILLER_0_1_613 ();
 sg13g2_fill_8 FILLER_0_1_621 ();
 sg13g2_fill_8 FILLER_0_1_629 ();
 sg13g2_fill_8 FILLER_0_1_637 ();
 sg13g2_fill_8 FILLER_0_1_645 ();
 sg13g2_fill_8 FILLER_0_1_653 ();
 sg13g2_fill_8 FILLER_0_1_661 ();
 sg13g2_fill_8 FILLER_0_1_669 ();
 sg13g2_fill_4 FILLER_0_1_677 ();
 sg13g2_fill_2 FILLER_0_1_681 ();
 sg13g2_fill_2 FILLER_0_1_709 ();
 sg13g2_fill_8 FILLER_0_1_716 ();
 sg13g2_fill_8 FILLER_0_1_724 ();
 sg13g2_fill_8 FILLER_0_1_732 ();
 sg13g2_fill_1 FILLER_0_1_740 ();
 sg13g2_fill_8 FILLER_0_1_767 ();
 sg13g2_fill_8 FILLER_0_1_775 ();
 sg13g2_fill_8 FILLER_0_1_783 ();
 sg13g2_fill_8 FILLER_0_1_791 ();
 sg13g2_fill_8 FILLER_0_1_799 ();
 sg13g2_fill_2 FILLER_0_1_807 ();
 sg13g2_fill_2 FILLER_0_1_835 ();
 sg13g2_fill_2 FILLER_0_1_842 ();
 sg13g2_fill_8 FILLER_0_1_848 ();
 sg13g2_fill_2 FILLER_0_1_856 ();
 sg13g2_fill_1 FILLER_0_1_858 ();
 sg13g2_fill_2 FILLER_0_1_864 ();
 sg13g2_fill_8 FILLER_0_1_892 ();
 sg13g2_fill_4 FILLER_0_1_900 ();
 sg13g2_fill_1 FILLER_0_1_904 ();
 sg13g2_fill_2 FILLER_0_1_909 ();
 sg13g2_fill_8 FILLER_0_1_937 ();
 sg13g2_fill_2 FILLER_0_1_945 ();
 sg13g2_fill_1 FILLER_0_1_947 ();
 sg13g2_fill_2 FILLER_0_1_953 ();
 sg13g2_fill_8 FILLER_0_1_959 ();
 sg13g2_fill_8 FILLER_0_1_967 ();
 sg13g2_fill_4 FILLER_0_1_975 ();
 sg13g2_fill_1 FILLER_0_1_979 ();
 sg13g2_fill_8 FILLER_0_1_1006 ();
 sg13g2_fill_2 FILLER_0_1_1014 ();
 sg13g2_fill_4 FILLER_0_1_1042 ();
 sg13g2_fill_1 FILLER_0_1_1046 ();
 sg13g2_fill_4 FILLER_0_1_1073 ();
 sg13g2_fill_1 FILLER_0_1_1077 ();
 sg13g2_fill_8 FILLER_0_1_1082 ();
 sg13g2_fill_8 FILLER_0_1_1093 ();
 sg13g2_fill_4 FILLER_0_1_1101 ();
 sg13g2_fill_2 FILLER_0_1_1105 ();
 sg13g2_fill_2 FILLER_0_1_1112 ();
 sg13g2_fill_2 FILLER_0_1_1118 ();
 sg13g2_fill_4 FILLER_0_1_1125 ();
 sg13g2_fill_8 FILLER_0_1_1155 ();
 sg13g2_fill_8 FILLER_0_1_1163 ();
 sg13g2_fill_8 FILLER_0_1_1171 ();
 sg13g2_fill_8 FILLER_0_1_1179 ();
 sg13g2_fill_8 FILLER_0_1_1187 ();
 sg13g2_fill_8 FILLER_0_1_1195 ();
 sg13g2_fill_8 FILLER_0_1_1203 ();
 sg13g2_fill_8 FILLER_0_1_1211 ();
 sg13g2_fill_8 FILLER_0_1_1219 ();
 sg13g2_fill_8 FILLER_0_1_1227 ();
 sg13g2_fill_8 FILLER_0_1_1235 ();
 sg13g2_fill_8 FILLER_0_1_1243 ();
 sg13g2_fill_8 FILLER_0_1_1251 ();
 sg13g2_fill_8 FILLER_0_1_1259 ();
 sg13g2_fill_8 FILLER_0_1_1267 ();
 sg13g2_fill_8 FILLER_0_1_1275 ();
 sg13g2_fill_8 FILLER_0_1_1283 ();
 sg13g2_fill_4 FILLER_0_1_1291 ();
 sg13g2_fill_2 FILLER_0_1_1295 ();
 sg13g2_fill_8 FILLER_0_2_0 ();
 sg13g2_fill_8 FILLER_0_2_8 ();
 sg13g2_fill_8 FILLER_0_2_16 ();
 sg13g2_fill_8 FILLER_0_2_24 ();
 sg13g2_fill_8 FILLER_0_2_32 ();
 sg13g2_fill_8 FILLER_0_2_40 ();
 sg13g2_fill_8 FILLER_0_2_48 ();
 sg13g2_fill_8 FILLER_0_2_56 ();
 sg13g2_fill_8 FILLER_0_2_64 ();
 sg13g2_fill_8 FILLER_0_2_72 ();
 sg13g2_fill_8 FILLER_0_2_80 ();
 sg13g2_fill_8 FILLER_0_2_88 ();
 sg13g2_fill_8 FILLER_0_2_96 ();
 sg13g2_fill_8 FILLER_0_2_104 ();
 sg13g2_fill_8 FILLER_0_2_112 ();
 sg13g2_fill_8 FILLER_0_2_120 ();
 sg13g2_fill_8 FILLER_0_2_128 ();
 sg13g2_fill_8 FILLER_0_2_136 ();
 sg13g2_fill_8 FILLER_0_2_144 ();
 sg13g2_fill_8 FILLER_0_2_152 ();
 sg13g2_fill_8 FILLER_0_2_160 ();
 sg13g2_fill_8 FILLER_0_2_168 ();
 sg13g2_fill_8 FILLER_0_2_176 ();
 sg13g2_fill_8 FILLER_0_2_184 ();
 sg13g2_fill_8 FILLER_0_2_192 ();
 sg13g2_fill_8 FILLER_0_2_200 ();
 sg13g2_fill_8 FILLER_0_2_208 ();
 sg13g2_fill_8 FILLER_0_2_216 ();
 sg13g2_fill_8 FILLER_0_2_224 ();
 sg13g2_fill_8 FILLER_0_2_232 ();
 sg13g2_fill_8 FILLER_0_2_240 ();
 sg13g2_fill_8 FILLER_0_2_248 ();
 sg13g2_fill_8 FILLER_0_2_256 ();
 sg13g2_fill_8 FILLER_0_2_264 ();
 sg13g2_fill_8 FILLER_0_2_272 ();
 sg13g2_fill_8 FILLER_0_2_280 ();
 sg13g2_fill_8 FILLER_0_2_288 ();
 sg13g2_fill_8 FILLER_0_2_296 ();
 sg13g2_fill_8 FILLER_0_2_304 ();
 sg13g2_fill_8 FILLER_0_2_312 ();
 sg13g2_fill_8 FILLER_0_2_320 ();
 sg13g2_fill_8 FILLER_0_2_328 ();
 sg13g2_fill_8 FILLER_0_2_336 ();
 sg13g2_fill_8 FILLER_0_2_344 ();
 sg13g2_fill_8 FILLER_0_2_352 ();
 sg13g2_fill_8 FILLER_0_2_360 ();
 sg13g2_fill_8 FILLER_0_2_368 ();
 sg13g2_fill_8 FILLER_0_2_376 ();
 sg13g2_fill_8 FILLER_0_2_384 ();
 sg13g2_fill_8 FILLER_0_2_392 ();
 sg13g2_fill_8 FILLER_0_2_400 ();
 sg13g2_fill_8 FILLER_0_2_408 ();
 sg13g2_fill_8 FILLER_0_2_416 ();
 sg13g2_fill_8 FILLER_0_2_424 ();
 sg13g2_fill_8 FILLER_0_2_432 ();
 sg13g2_fill_8 FILLER_0_2_440 ();
 sg13g2_fill_8 FILLER_0_2_448 ();
 sg13g2_fill_8 FILLER_0_2_456 ();
 sg13g2_fill_8 FILLER_0_2_464 ();
 sg13g2_fill_8 FILLER_0_2_472 ();
 sg13g2_fill_8 FILLER_0_2_480 ();
 sg13g2_fill_8 FILLER_0_2_488 ();
 sg13g2_fill_8 FILLER_0_2_496 ();
 sg13g2_fill_8 FILLER_0_2_504 ();
 sg13g2_fill_8 FILLER_0_2_512 ();
 sg13g2_fill_8 FILLER_0_2_520 ();
 sg13g2_fill_8 FILLER_0_2_528 ();
 sg13g2_fill_8 FILLER_0_2_536 ();
 sg13g2_fill_2 FILLER_0_2_549 ();
 sg13g2_fill_2 FILLER_0_2_577 ();
 sg13g2_fill_2 FILLER_0_2_583 ();
 sg13g2_fill_2 FILLER_0_2_590 ();
 sg13g2_fill_8 FILLER_0_2_618 ();
 sg13g2_fill_8 FILLER_0_2_626 ();
 sg13g2_fill_8 FILLER_0_2_634 ();
 sg13g2_fill_8 FILLER_0_2_642 ();
 sg13g2_fill_8 FILLER_0_2_650 ();
 sg13g2_fill_4 FILLER_0_2_658 ();
 sg13g2_fill_2 FILLER_0_2_662 ();
 sg13g2_fill_1 FILLER_0_2_664 ();
 sg13g2_fill_2 FILLER_0_2_691 ();
 sg13g2_fill_4 FILLER_0_2_697 ();
 sg13g2_fill_4 FILLER_0_2_727 ();
 sg13g2_fill_2 FILLER_0_2_757 ();
 sg13g2_fill_8 FILLER_0_2_764 ();
 sg13g2_fill_8 FILLER_0_2_772 ();
 sg13g2_fill_4 FILLER_0_2_780 ();
 sg13g2_fill_2 FILLER_0_2_810 ();
 sg13g2_fill_2 FILLER_0_2_817 ();
 sg13g2_fill_1 FILLER_0_2_819 ();
 sg13g2_fill_4 FILLER_0_2_824 ();
 sg13g2_fill_1 FILLER_0_2_828 ();
 sg13g2_fill_4 FILLER_0_2_855 ();
 sg13g2_fill_1 FILLER_0_2_859 ();
 sg13g2_fill_4 FILLER_0_2_886 ();
 sg13g2_fill_1 FILLER_0_2_890 ();
 sg13g2_fill_4 FILLER_0_2_895 ();
 sg13g2_fill_2 FILLER_0_2_899 ();
 sg13g2_fill_1 FILLER_0_2_901 ();
 sg13g2_fill_2 FILLER_0_2_928 ();
 sg13g2_fill_8 FILLER_0_2_934 ();
 sg13g2_fill_2 FILLER_0_2_942 ();
 sg13g2_fill_4 FILLER_0_2_970 ();
 sg13g2_fill_2 FILLER_0_2_974 ();
 sg13g2_fill_1 FILLER_0_2_976 ();
 sg13g2_fill_2 FILLER_0_2_998 ();
 sg13g2_fill_8 FILLER_0_2_1005 ();
 sg13g2_fill_2 FILLER_0_2_1018 ();
 sg13g2_fill_8 FILLER_0_2_1024 ();
 sg13g2_fill_8 FILLER_0_2_1032 ();
 sg13g2_fill_8 FILLER_0_2_1040 ();
 sg13g2_fill_8 FILLER_0_2_1048 ();
 sg13g2_fill_8 FILLER_0_2_1056 ();
 sg13g2_fill_2 FILLER_0_2_1069 ();
 sg13g2_fill_8 FILLER_0_2_1097 ();
 sg13g2_fill_1 FILLER_0_2_1105 ();
 sg13g2_fill_4 FILLER_0_2_1132 ();
 sg13g2_fill_8 FILLER_0_2_1157 ();
 sg13g2_fill_8 FILLER_0_2_1165 ();
 sg13g2_fill_8 FILLER_0_2_1173 ();
 sg13g2_fill_8 FILLER_0_2_1181 ();
 sg13g2_fill_8 FILLER_0_2_1189 ();
 sg13g2_fill_8 FILLER_0_2_1197 ();
 sg13g2_fill_8 FILLER_0_2_1205 ();
 sg13g2_fill_8 FILLER_0_2_1213 ();
 sg13g2_fill_8 FILLER_0_2_1221 ();
 sg13g2_fill_8 FILLER_0_2_1229 ();
 sg13g2_fill_8 FILLER_0_2_1237 ();
 sg13g2_fill_8 FILLER_0_2_1245 ();
 sg13g2_fill_8 FILLER_0_2_1253 ();
 sg13g2_fill_8 FILLER_0_2_1261 ();
 sg13g2_fill_8 FILLER_0_2_1269 ();
 sg13g2_fill_8 FILLER_0_2_1277 ();
 sg13g2_fill_8 FILLER_0_2_1285 ();
 sg13g2_fill_4 FILLER_0_2_1293 ();
 sg13g2_fill_8 FILLER_0_3_0 ();
 sg13g2_fill_8 FILLER_0_3_8 ();
 sg13g2_fill_8 FILLER_0_3_16 ();
 sg13g2_fill_8 FILLER_0_3_24 ();
 sg13g2_fill_8 FILLER_0_3_32 ();
 sg13g2_fill_8 FILLER_0_3_40 ();
 sg13g2_fill_8 FILLER_0_3_48 ();
 sg13g2_fill_8 FILLER_0_3_56 ();
 sg13g2_fill_8 FILLER_0_3_64 ();
 sg13g2_fill_8 FILLER_0_3_72 ();
 sg13g2_fill_8 FILLER_0_3_80 ();
 sg13g2_fill_8 FILLER_0_3_88 ();
 sg13g2_fill_8 FILLER_0_3_96 ();
 sg13g2_fill_8 FILLER_0_3_104 ();
 sg13g2_fill_8 FILLER_0_3_112 ();
 sg13g2_fill_8 FILLER_0_3_120 ();
 sg13g2_fill_8 FILLER_0_3_128 ();
 sg13g2_fill_8 FILLER_0_3_136 ();
 sg13g2_fill_8 FILLER_0_3_144 ();
 sg13g2_fill_8 FILLER_0_3_152 ();
 sg13g2_fill_8 FILLER_0_3_160 ();
 sg13g2_fill_8 FILLER_0_3_168 ();
 sg13g2_fill_8 FILLER_0_3_176 ();
 sg13g2_fill_8 FILLER_0_3_184 ();
 sg13g2_fill_8 FILLER_0_3_192 ();
 sg13g2_fill_8 FILLER_0_3_200 ();
 sg13g2_fill_8 FILLER_0_3_208 ();
 sg13g2_fill_8 FILLER_0_3_216 ();
 sg13g2_fill_8 FILLER_0_3_224 ();
 sg13g2_fill_8 FILLER_0_3_232 ();
 sg13g2_fill_8 FILLER_0_3_240 ();
 sg13g2_fill_8 FILLER_0_3_248 ();
 sg13g2_fill_8 FILLER_0_3_256 ();
 sg13g2_fill_8 FILLER_0_3_264 ();
 sg13g2_fill_8 FILLER_0_3_272 ();
 sg13g2_fill_8 FILLER_0_3_280 ();
 sg13g2_fill_8 FILLER_0_3_288 ();
 sg13g2_fill_8 FILLER_0_3_296 ();
 sg13g2_fill_8 FILLER_0_3_304 ();
 sg13g2_fill_8 FILLER_0_3_312 ();
 sg13g2_fill_8 FILLER_0_3_320 ();
 sg13g2_fill_8 FILLER_0_3_328 ();
 sg13g2_fill_8 FILLER_0_3_336 ();
 sg13g2_fill_8 FILLER_0_3_344 ();
 sg13g2_fill_8 FILLER_0_3_352 ();
 sg13g2_fill_8 FILLER_0_3_360 ();
 sg13g2_fill_8 FILLER_0_3_368 ();
 sg13g2_fill_8 FILLER_0_3_376 ();
 sg13g2_fill_8 FILLER_0_3_384 ();
 sg13g2_fill_8 FILLER_0_3_392 ();
 sg13g2_fill_8 FILLER_0_3_400 ();
 sg13g2_fill_8 FILLER_0_3_408 ();
 sg13g2_fill_8 FILLER_0_3_416 ();
 sg13g2_fill_8 FILLER_0_3_424 ();
 sg13g2_fill_8 FILLER_0_3_432 ();
 sg13g2_fill_8 FILLER_0_3_440 ();
 sg13g2_fill_8 FILLER_0_3_448 ();
 sg13g2_fill_8 FILLER_0_3_456 ();
 sg13g2_fill_8 FILLER_0_3_464 ();
 sg13g2_fill_8 FILLER_0_3_472 ();
 sg13g2_fill_8 FILLER_0_3_480 ();
 sg13g2_fill_8 FILLER_0_3_488 ();
 sg13g2_fill_8 FILLER_0_3_496 ();
 sg13g2_fill_8 FILLER_0_3_504 ();
 sg13g2_fill_8 FILLER_0_3_512 ();
 sg13g2_fill_8 FILLER_0_3_520 ();
 sg13g2_fill_8 FILLER_0_3_528 ();
 sg13g2_fill_8 FILLER_0_3_536 ();
 sg13g2_fill_8 FILLER_0_3_544 ();
 sg13g2_fill_1 FILLER_0_3_552 ();
 sg13g2_fill_2 FILLER_0_3_558 ();
 sg13g2_fill_2 FILLER_0_3_564 ();
 sg13g2_fill_1 FILLER_0_3_566 ();
 sg13g2_fill_2 FILLER_0_3_588 ();
 sg13g2_fill_4 FILLER_0_3_594 ();
 sg13g2_fill_1 FILLER_0_3_598 ();
 sg13g2_fill_8 FILLER_0_3_620 ();
 sg13g2_fill_8 FILLER_0_3_628 ();
 sg13g2_fill_2 FILLER_0_3_636 ();
 sg13g2_fill_2 FILLER_0_3_643 ();
 sg13g2_fill_1 FILLER_0_3_645 ();
 sg13g2_fill_2 FILLER_0_3_651 ();
 sg13g2_fill_2 FILLER_0_3_679 ();
 sg13g2_fill_2 FILLER_0_3_685 ();
 sg13g2_fill_1 FILLER_0_3_687 ();
 sg13g2_fill_4 FILLER_0_3_693 ();
 sg13g2_fill_2 FILLER_0_3_697 ();
 sg13g2_fill_8 FILLER_0_3_720 ();
 sg13g2_fill_1 FILLER_0_3_728 ();
 sg13g2_fill_4 FILLER_0_3_734 ();
 sg13g2_fill_8 FILLER_0_3_742 ();
 sg13g2_fill_8 FILLER_0_3_750 ();
 sg13g2_fill_8 FILLER_0_3_762 ();
 sg13g2_fill_8 FILLER_0_3_770 ();
 sg13g2_fill_8 FILLER_0_3_778 ();
 sg13g2_fill_4 FILLER_0_3_786 ();
 sg13g2_fill_2 FILLER_0_3_790 ();
 sg13g2_fill_1 FILLER_0_3_792 ();
 sg13g2_fill_4 FILLER_0_3_797 ();
 sg13g2_fill_2 FILLER_0_3_806 ();
 sg13g2_fill_2 FILLER_0_3_834 ();
 sg13g2_fill_1 FILLER_0_3_836 ();
 sg13g2_fill_8 FILLER_0_3_858 ();
 sg13g2_fill_2 FILLER_0_3_866 ();
 sg13g2_fill_1 FILLER_0_3_868 ();
 sg13g2_fill_2 FILLER_0_3_873 ();
 sg13g2_fill_2 FILLER_0_3_880 ();
 sg13g2_fill_4 FILLER_0_3_892 ();
 sg13g2_fill_2 FILLER_0_3_896 ();
 sg13g2_fill_1 FILLER_0_3_898 ();
 sg13g2_fill_8 FILLER_0_3_904 ();
 sg13g2_fill_1 FILLER_0_3_912 ();
 sg13g2_fill_2 FILLER_0_3_918 ();
 sg13g2_fill_2 FILLER_0_3_925 ();
 sg13g2_fill_1 FILLER_0_3_927 ();
 sg13g2_fill_8 FILLER_0_3_934 ();
 sg13g2_fill_2 FILLER_0_3_942 ();
 sg13g2_fill_2 FILLER_0_3_970 ();
 sg13g2_fill_2 FILLER_0_3_998 ();
 sg13g2_fill_8 FILLER_0_3_1004 ();
 sg13g2_fill_4 FILLER_0_3_1012 ();
 sg13g2_fill_1 FILLER_0_3_1016 ();
 sg13g2_fill_8 FILLER_0_3_1023 ();
 sg13g2_fill_8 FILLER_0_3_1031 ();
 sg13g2_fill_8 FILLER_0_3_1039 ();
 sg13g2_fill_2 FILLER_0_3_1047 ();
 sg13g2_fill_1 FILLER_0_3_1049 ();
 sg13g2_fill_8 FILLER_0_3_1055 ();
 sg13g2_fill_1 FILLER_0_3_1063 ();
 sg13g2_fill_2 FILLER_0_3_1068 ();
 sg13g2_fill_8 FILLER_0_3_1074 ();
 sg13g2_fill_8 FILLER_0_3_1082 ();
 sg13g2_fill_8 FILLER_0_3_1090 ();
 sg13g2_fill_1 FILLER_0_3_1098 ();
 sg13g2_fill_8 FILLER_0_3_1103 ();
 sg13g2_fill_2 FILLER_0_3_1111 ();
 sg13g2_fill_1 FILLER_0_3_1113 ();
 sg13g2_fill_2 FILLER_0_3_1117 ();
 sg13g2_fill_8 FILLER_0_3_1123 ();
 sg13g2_fill_8 FILLER_0_3_1152 ();
 sg13g2_fill_8 FILLER_0_3_1160 ();
 sg13g2_fill_8 FILLER_0_3_1168 ();
 sg13g2_fill_8 FILLER_0_3_1176 ();
 sg13g2_fill_8 FILLER_0_3_1184 ();
 sg13g2_fill_8 FILLER_0_3_1192 ();
 sg13g2_fill_8 FILLER_0_3_1200 ();
 sg13g2_fill_8 FILLER_0_3_1208 ();
 sg13g2_fill_8 FILLER_0_3_1216 ();
 sg13g2_fill_8 FILLER_0_3_1224 ();
 sg13g2_fill_8 FILLER_0_3_1232 ();
 sg13g2_fill_8 FILLER_0_3_1240 ();
 sg13g2_fill_8 FILLER_0_3_1248 ();
 sg13g2_fill_8 FILLER_0_3_1256 ();
 sg13g2_fill_8 FILLER_0_3_1264 ();
 sg13g2_fill_8 FILLER_0_3_1272 ();
 sg13g2_fill_8 FILLER_0_3_1280 ();
 sg13g2_fill_8 FILLER_0_3_1288 ();
 sg13g2_fill_1 FILLER_0_3_1296 ();
 sg13g2_fill_8 FILLER_0_4_0 ();
 sg13g2_fill_8 FILLER_0_4_8 ();
 sg13g2_fill_8 FILLER_0_4_16 ();
 sg13g2_fill_8 FILLER_0_4_24 ();
 sg13g2_fill_8 FILLER_0_4_32 ();
 sg13g2_fill_8 FILLER_0_4_40 ();
 sg13g2_fill_8 FILLER_0_4_48 ();
 sg13g2_fill_8 FILLER_0_4_56 ();
 sg13g2_fill_8 FILLER_0_4_64 ();
 sg13g2_fill_8 FILLER_0_4_72 ();
 sg13g2_fill_8 FILLER_0_4_80 ();
 sg13g2_fill_8 FILLER_0_4_88 ();
 sg13g2_fill_8 FILLER_0_4_96 ();
 sg13g2_fill_8 FILLER_0_4_104 ();
 sg13g2_fill_8 FILLER_0_4_112 ();
 sg13g2_fill_8 FILLER_0_4_120 ();
 sg13g2_fill_8 FILLER_0_4_128 ();
 sg13g2_fill_8 FILLER_0_4_136 ();
 sg13g2_fill_8 FILLER_0_4_144 ();
 sg13g2_fill_8 FILLER_0_4_152 ();
 sg13g2_fill_8 FILLER_0_4_160 ();
 sg13g2_fill_8 FILLER_0_4_168 ();
 sg13g2_fill_8 FILLER_0_4_176 ();
 sg13g2_fill_8 FILLER_0_4_184 ();
 sg13g2_fill_8 FILLER_0_4_192 ();
 sg13g2_fill_8 FILLER_0_4_200 ();
 sg13g2_fill_8 FILLER_0_4_208 ();
 sg13g2_fill_8 FILLER_0_4_216 ();
 sg13g2_fill_8 FILLER_0_4_224 ();
 sg13g2_fill_8 FILLER_0_4_232 ();
 sg13g2_fill_8 FILLER_0_4_240 ();
 sg13g2_fill_8 FILLER_0_4_248 ();
 sg13g2_fill_8 FILLER_0_4_256 ();
 sg13g2_fill_8 FILLER_0_4_264 ();
 sg13g2_fill_8 FILLER_0_4_272 ();
 sg13g2_fill_8 FILLER_0_4_280 ();
 sg13g2_fill_8 FILLER_0_4_288 ();
 sg13g2_fill_8 FILLER_0_4_296 ();
 sg13g2_fill_8 FILLER_0_4_304 ();
 sg13g2_fill_8 FILLER_0_4_312 ();
 sg13g2_fill_8 FILLER_0_4_320 ();
 sg13g2_fill_8 FILLER_0_4_328 ();
 sg13g2_fill_8 FILLER_0_4_336 ();
 sg13g2_fill_8 FILLER_0_4_344 ();
 sg13g2_fill_8 FILLER_0_4_352 ();
 sg13g2_fill_8 FILLER_0_4_360 ();
 sg13g2_fill_8 FILLER_0_4_368 ();
 sg13g2_fill_8 FILLER_0_4_376 ();
 sg13g2_fill_8 FILLER_0_4_384 ();
 sg13g2_fill_8 FILLER_0_4_392 ();
 sg13g2_fill_8 FILLER_0_4_400 ();
 sg13g2_fill_8 FILLER_0_4_408 ();
 sg13g2_fill_8 FILLER_0_4_416 ();
 sg13g2_fill_8 FILLER_0_4_424 ();
 sg13g2_fill_8 FILLER_0_4_432 ();
 sg13g2_fill_8 FILLER_0_4_440 ();
 sg13g2_fill_8 FILLER_0_4_448 ();
 sg13g2_fill_8 FILLER_0_4_456 ();
 sg13g2_fill_8 FILLER_0_4_464 ();
 sg13g2_fill_8 FILLER_0_4_472 ();
 sg13g2_fill_8 FILLER_0_4_480 ();
 sg13g2_fill_8 FILLER_0_4_488 ();
 sg13g2_fill_8 FILLER_0_4_496 ();
 sg13g2_fill_8 FILLER_0_4_504 ();
 sg13g2_fill_8 FILLER_0_4_512 ();
 sg13g2_fill_8 FILLER_0_4_520 ();
 sg13g2_fill_8 FILLER_0_4_528 ();
 sg13g2_fill_8 FILLER_0_4_536 ();
 sg13g2_fill_8 FILLER_0_4_544 ();
 sg13g2_fill_8 FILLER_0_4_552 ();
 sg13g2_fill_8 FILLER_0_4_560 ();
 sg13g2_fill_8 FILLER_0_4_568 ();
 sg13g2_fill_8 FILLER_0_4_576 ();
 sg13g2_fill_4 FILLER_0_4_584 ();
 sg13g2_fill_8 FILLER_0_4_593 ();
 sg13g2_fill_8 FILLER_0_4_601 ();
 sg13g2_fill_8 FILLER_0_4_609 ();
 sg13g2_fill_8 FILLER_0_4_617 ();
 sg13g2_fill_8 FILLER_0_4_625 ();
 sg13g2_fill_8 FILLER_0_4_633 ();
 sg13g2_fill_8 FILLER_0_4_641 ();
 sg13g2_fill_2 FILLER_0_4_649 ();
 sg13g2_fill_1 FILLER_0_4_651 ();
 sg13g2_fill_8 FILLER_0_4_656 ();
 sg13g2_fill_8 FILLER_0_4_664 ();
 sg13g2_fill_2 FILLER_0_4_677 ();
 sg13g2_fill_8 FILLER_0_4_689 ();
 sg13g2_fill_8 FILLER_0_4_697 ();
 sg13g2_fill_4 FILLER_0_4_705 ();
 sg13g2_fill_8 FILLER_0_4_715 ();
 sg13g2_fill_8 FILLER_0_4_723 ();
 sg13g2_fill_8 FILLER_0_4_731 ();
 sg13g2_fill_8 FILLER_0_4_739 ();
 sg13g2_fill_1 FILLER_0_4_747 ();
 sg13g2_fill_8 FILLER_0_4_758 ();
 sg13g2_fill_8 FILLER_0_4_766 ();
 sg13g2_fill_8 FILLER_0_4_774 ();
 sg13g2_fill_8 FILLER_0_4_782 ();
 sg13g2_fill_2 FILLER_0_4_790 ();
 sg13g2_fill_1 FILLER_0_4_792 ();
 sg13g2_fill_2 FILLER_0_4_798 ();
 sg13g2_fill_8 FILLER_0_4_804 ();
 sg13g2_fill_8 FILLER_0_4_812 ();
 sg13g2_fill_2 FILLER_0_4_820 ();
 sg13g2_fill_1 FILLER_0_4_822 ();
 sg13g2_fill_8 FILLER_0_4_844 ();
 sg13g2_fill_8 FILLER_0_4_852 ();
 sg13g2_fill_8 FILLER_0_4_860 ();
 sg13g2_fill_8 FILLER_0_4_868 ();
 sg13g2_fill_8 FILLER_0_4_876 ();
 sg13g2_fill_8 FILLER_0_4_884 ();
 sg13g2_fill_8 FILLER_0_4_892 ();
 sg13g2_fill_8 FILLER_0_4_900 ();
 sg13g2_fill_8 FILLER_0_4_908 ();
 sg13g2_fill_8 FILLER_0_4_916 ();
 sg13g2_fill_8 FILLER_0_4_924 ();
 sg13g2_fill_8 FILLER_0_4_932 ();
 sg13g2_fill_8 FILLER_0_4_940 ();
 sg13g2_fill_4 FILLER_0_4_953 ();
 sg13g2_fill_1 FILLER_0_4_957 ();
 sg13g2_fill_8 FILLER_0_4_962 ();
 sg13g2_fill_2 FILLER_0_4_975 ();
 sg13g2_fill_2 FILLER_0_4_998 ();
 sg13g2_fill_4 FILLER_0_4_1004 ();
 sg13g2_fill_2 FILLER_0_4_1008 ();
 sg13g2_fill_1 FILLER_0_4_1010 ();
 sg13g2_fill_2 FILLER_0_4_1016 ();
 sg13g2_fill_4 FILLER_0_4_1022 ();
 sg13g2_fill_2 FILLER_0_4_1026 ();
 sg13g2_fill_8 FILLER_0_4_1033 ();
 sg13g2_fill_2 FILLER_0_4_1041 ();
 sg13g2_fill_1 FILLER_0_4_1043 ();
 sg13g2_fill_2 FILLER_0_4_1070 ();
 sg13g2_fill_4 FILLER_0_4_1093 ();
 sg13g2_fill_2 FILLER_0_4_1097 ();
 sg13g2_fill_2 FILLER_0_4_1104 ();
 sg13g2_fill_2 FILLER_0_4_1132 ();
 sg13g2_fill_1 FILLER_0_4_1134 ();
 sg13g2_fill_2 FILLER_0_4_1139 ();
 sg13g2_fill_2 FILLER_0_4_1146 ();
 sg13g2_fill_8 FILLER_0_4_1174 ();
 sg13g2_fill_8 FILLER_0_4_1182 ();
 sg13g2_fill_8 FILLER_0_4_1190 ();
 sg13g2_fill_8 FILLER_0_4_1198 ();
 sg13g2_fill_8 FILLER_0_4_1206 ();
 sg13g2_fill_8 FILLER_0_4_1214 ();
 sg13g2_fill_8 FILLER_0_4_1222 ();
 sg13g2_fill_8 FILLER_0_4_1230 ();
 sg13g2_fill_8 FILLER_0_4_1238 ();
 sg13g2_fill_8 FILLER_0_4_1246 ();
 sg13g2_fill_8 FILLER_0_4_1254 ();
 sg13g2_fill_8 FILLER_0_4_1262 ();
 sg13g2_fill_8 FILLER_0_4_1270 ();
 sg13g2_fill_8 FILLER_0_4_1278 ();
 sg13g2_fill_8 FILLER_0_4_1286 ();
 sg13g2_fill_2 FILLER_0_4_1294 ();
 sg13g2_fill_1 FILLER_0_4_1296 ();
 sg13g2_fill_8 FILLER_0_5_0 ();
 sg13g2_fill_8 FILLER_0_5_8 ();
 sg13g2_fill_8 FILLER_0_5_16 ();
 sg13g2_fill_8 FILLER_0_5_24 ();
 sg13g2_fill_8 FILLER_0_5_32 ();
 sg13g2_fill_8 FILLER_0_5_40 ();
 sg13g2_fill_8 FILLER_0_5_48 ();
 sg13g2_fill_8 FILLER_0_5_56 ();
 sg13g2_fill_8 FILLER_0_5_64 ();
 sg13g2_fill_8 FILLER_0_5_72 ();
 sg13g2_fill_8 FILLER_0_5_80 ();
 sg13g2_fill_8 FILLER_0_5_88 ();
 sg13g2_fill_8 FILLER_0_5_96 ();
 sg13g2_fill_8 FILLER_0_5_104 ();
 sg13g2_fill_8 FILLER_0_5_112 ();
 sg13g2_fill_8 FILLER_0_5_120 ();
 sg13g2_fill_8 FILLER_0_5_128 ();
 sg13g2_fill_8 FILLER_0_5_136 ();
 sg13g2_fill_8 FILLER_0_5_144 ();
 sg13g2_fill_8 FILLER_0_5_152 ();
 sg13g2_fill_8 FILLER_0_5_160 ();
 sg13g2_fill_8 FILLER_0_5_168 ();
 sg13g2_fill_8 FILLER_0_5_176 ();
 sg13g2_fill_8 FILLER_0_5_184 ();
 sg13g2_fill_8 FILLER_0_5_192 ();
 sg13g2_fill_8 FILLER_0_5_200 ();
 sg13g2_fill_8 FILLER_0_5_208 ();
 sg13g2_fill_8 FILLER_0_5_216 ();
 sg13g2_fill_8 FILLER_0_5_224 ();
 sg13g2_fill_8 FILLER_0_5_232 ();
 sg13g2_fill_8 FILLER_0_5_240 ();
 sg13g2_fill_8 FILLER_0_5_248 ();
 sg13g2_fill_8 FILLER_0_5_256 ();
 sg13g2_fill_8 FILLER_0_5_264 ();
 sg13g2_fill_8 FILLER_0_5_272 ();
 sg13g2_fill_8 FILLER_0_5_280 ();
 sg13g2_fill_8 FILLER_0_5_288 ();
 sg13g2_fill_8 FILLER_0_5_296 ();
 sg13g2_fill_8 FILLER_0_5_304 ();
 sg13g2_fill_8 FILLER_0_5_312 ();
 sg13g2_fill_8 FILLER_0_5_320 ();
 sg13g2_fill_8 FILLER_0_5_328 ();
 sg13g2_fill_8 FILLER_0_5_336 ();
 sg13g2_fill_8 FILLER_0_5_344 ();
 sg13g2_fill_4 FILLER_0_5_352 ();
 sg13g2_fill_2 FILLER_0_5_356 ();
 sg13g2_fill_8 FILLER_0_5_362 ();
 sg13g2_fill_8 FILLER_0_5_370 ();
 sg13g2_fill_8 FILLER_0_5_378 ();
 sg13g2_fill_8 FILLER_0_5_386 ();
 sg13g2_fill_8 FILLER_0_5_394 ();
 sg13g2_fill_4 FILLER_0_5_402 ();
 sg13g2_fill_2 FILLER_0_5_406 ();
 sg13g2_fill_8 FILLER_0_5_434 ();
 sg13g2_fill_8 FILLER_0_5_442 ();
 sg13g2_fill_8 FILLER_0_5_450 ();
 sg13g2_fill_8 FILLER_0_5_458 ();
 sg13g2_fill_2 FILLER_0_5_466 ();
 sg13g2_fill_8 FILLER_0_5_473 ();
 sg13g2_fill_8 FILLER_0_5_481 ();
 sg13g2_fill_8 FILLER_0_5_489 ();
 sg13g2_fill_4 FILLER_0_5_497 ();
 sg13g2_fill_2 FILLER_0_5_501 ();
 sg13g2_fill_1 FILLER_0_5_503 ();
 sg13g2_fill_2 FILLER_0_5_530 ();
 sg13g2_fill_8 FILLER_0_5_537 ();
 sg13g2_fill_2 FILLER_0_5_545 ();
 sg13g2_fill_1 FILLER_0_5_547 ();
 sg13g2_fill_8 FILLER_0_5_553 ();
 sg13g2_fill_8 FILLER_0_5_561 ();
 sg13g2_fill_8 FILLER_0_5_569 ();
 sg13g2_fill_8 FILLER_0_5_577 ();
 sg13g2_fill_8 FILLER_0_5_585 ();
 sg13g2_fill_8 FILLER_0_5_593 ();
 sg13g2_fill_4 FILLER_0_5_601 ();
 sg13g2_fill_2 FILLER_0_5_605 ();
 sg13g2_fill_1 FILLER_0_5_607 ();
 sg13g2_fill_2 FILLER_0_5_613 ();
 sg13g2_fill_2 FILLER_0_5_619 ();
 sg13g2_fill_8 FILLER_0_5_647 ();
 sg13g2_fill_8 FILLER_0_5_655 ();
 sg13g2_fill_8 FILLER_0_5_663 ();
 sg13g2_fill_8 FILLER_0_5_671 ();
 sg13g2_fill_8 FILLER_0_5_679 ();
 sg13g2_fill_8 FILLER_0_5_687 ();
 sg13g2_fill_8 FILLER_0_5_695 ();
 sg13g2_fill_8 FILLER_0_5_703 ();
 sg13g2_fill_8 FILLER_0_5_711 ();
 sg13g2_fill_8 FILLER_0_5_719 ();
 sg13g2_fill_8 FILLER_0_5_727 ();
 sg13g2_fill_8 FILLER_0_5_735 ();
 sg13g2_fill_2 FILLER_0_5_743 ();
 sg13g2_fill_1 FILLER_0_5_745 ();
 sg13g2_fill_8 FILLER_0_5_767 ();
 sg13g2_fill_8 FILLER_0_5_775 ();
 sg13g2_fill_8 FILLER_0_5_783 ();
 sg13g2_fill_8 FILLER_0_5_791 ();
 sg13g2_fill_8 FILLER_0_5_799 ();
 sg13g2_fill_8 FILLER_0_5_807 ();
 sg13g2_fill_8 FILLER_0_5_815 ();
 sg13g2_fill_8 FILLER_0_5_823 ();
 sg13g2_fill_8 FILLER_0_5_831 ();
 sg13g2_fill_8 FILLER_0_5_839 ();
 sg13g2_fill_8 FILLER_0_5_847 ();
 sg13g2_fill_8 FILLER_0_5_855 ();
 sg13g2_fill_8 FILLER_0_5_863 ();
 sg13g2_fill_4 FILLER_0_5_871 ();
 sg13g2_fill_2 FILLER_0_5_875 ();
 sg13g2_fill_1 FILLER_0_5_877 ();
 sg13g2_fill_8 FILLER_0_5_899 ();
 sg13g2_fill_8 FILLER_0_5_907 ();
 sg13g2_fill_4 FILLER_0_5_915 ();
 sg13g2_fill_2 FILLER_0_5_919 ();
 sg13g2_fill_2 FILLER_0_5_942 ();
 sg13g2_fill_8 FILLER_0_5_949 ();
 sg13g2_fill_8 FILLER_0_5_957 ();
 sg13g2_fill_8 FILLER_0_5_965 ();
 sg13g2_fill_8 FILLER_0_5_973 ();
 sg13g2_fill_8 FILLER_0_5_981 ();
 sg13g2_fill_8 FILLER_0_5_989 ();
 sg13g2_fill_8 FILLER_0_5_997 ();
 sg13g2_fill_4 FILLER_0_5_1005 ();
 sg13g2_fill_2 FILLER_0_5_1009 ();
 sg13g2_fill_1 FILLER_0_5_1011 ();
 sg13g2_fill_8 FILLER_0_5_1038 ();
 sg13g2_fill_1 FILLER_0_5_1046 ();
 sg13g2_fill_4 FILLER_0_5_1052 ();
 sg13g2_fill_1 FILLER_0_5_1056 ();
 sg13g2_fill_2 FILLER_0_5_1062 ();
 sg13g2_fill_4 FILLER_0_5_1068 ();
 sg13g2_fill_1 FILLER_0_5_1072 ();
 sg13g2_fill_8 FILLER_0_5_1094 ();
 sg13g2_fill_8 FILLER_0_5_1102 ();
 sg13g2_fill_8 FILLER_0_5_1110 ();
 sg13g2_fill_8 FILLER_0_5_1118 ();
 sg13g2_fill_8 FILLER_0_5_1126 ();
 sg13g2_fill_8 FILLER_0_5_1134 ();
 sg13g2_fill_8 FILLER_0_5_1142 ();
 sg13g2_fill_8 FILLER_0_5_1150 ();
 sg13g2_fill_8 FILLER_0_5_1158 ();
 sg13g2_fill_8 FILLER_0_5_1166 ();
 sg13g2_fill_2 FILLER_0_5_1174 ();
 sg13g2_fill_8 FILLER_0_5_1202 ();
 sg13g2_fill_8 FILLER_0_5_1210 ();
 sg13g2_fill_8 FILLER_0_5_1218 ();
 sg13g2_fill_8 FILLER_0_5_1226 ();
 sg13g2_fill_8 FILLER_0_5_1234 ();
 sg13g2_fill_8 FILLER_0_5_1242 ();
 sg13g2_fill_8 FILLER_0_5_1250 ();
 sg13g2_fill_8 FILLER_0_5_1258 ();
 sg13g2_fill_8 FILLER_0_5_1266 ();
 sg13g2_fill_8 FILLER_0_5_1274 ();
 sg13g2_fill_8 FILLER_0_5_1282 ();
 sg13g2_fill_4 FILLER_0_5_1290 ();
 sg13g2_fill_2 FILLER_0_5_1294 ();
 sg13g2_fill_1 FILLER_0_5_1296 ();
 sg13g2_fill_8 FILLER_0_6_0 ();
 sg13g2_fill_8 FILLER_0_6_8 ();
 sg13g2_fill_8 FILLER_0_6_16 ();
 sg13g2_fill_8 FILLER_0_6_24 ();
 sg13g2_fill_8 FILLER_0_6_32 ();
 sg13g2_fill_8 FILLER_0_6_40 ();
 sg13g2_fill_8 FILLER_0_6_48 ();
 sg13g2_fill_8 FILLER_0_6_56 ();
 sg13g2_fill_8 FILLER_0_6_64 ();
 sg13g2_fill_8 FILLER_0_6_72 ();
 sg13g2_fill_8 FILLER_0_6_80 ();
 sg13g2_fill_8 FILLER_0_6_88 ();
 sg13g2_fill_8 FILLER_0_6_96 ();
 sg13g2_fill_8 FILLER_0_6_104 ();
 sg13g2_fill_8 FILLER_0_6_112 ();
 sg13g2_fill_8 FILLER_0_6_120 ();
 sg13g2_fill_8 FILLER_0_6_128 ();
 sg13g2_fill_8 FILLER_0_6_136 ();
 sg13g2_fill_8 FILLER_0_6_144 ();
 sg13g2_fill_8 FILLER_0_6_152 ();
 sg13g2_fill_8 FILLER_0_6_160 ();
 sg13g2_fill_8 FILLER_0_6_168 ();
 sg13g2_fill_8 FILLER_0_6_176 ();
 sg13g2_fill_8 FILLER_0_6_184 ();
 sg13g2_fill_8 FILLER_0_6_192 ();
 sg13g2_fill_8 FILLER_0_6_200 ();
 sg13g2_fill_8 FILLER_0_6_208 ();
 sg13g2_fill_8 FILLER_0_6_216 ();
 sg13g2_fill_8 FILLER_0_6_224 ();
 sg13g2_fill_8 FILLER_0_6_232 ();
 sg13g2_fill_8 FILLER_0_6_240 ();
 sg13g2_fill_8 FILLER_0_6_248 ();
 sg13g2_fill_8 FILLER_0_6_256 ();
 sg13g2_fill_8 FILLER_0_6_264 ();
 sg13g2_fill_8 FILLER_0_6_272 ();
 sg13g2_fill_8 FILLER_0_6_280 ();
 sg13g2_fill_8 FILLER_0_6_288 ();
 sg13g2_fill_8 FILLER_0_6_296 ();
 sg13g2_fill_8 FILLER_0_6_304 ();
 sg13g2_fill_8 FILLER_0_6_312 ();
 sg13g2_fill_8 FILLER_0_6_320 ();
 sg13g2_fill_8 FILLER_0_6_328 ();
 sg13g2_fill_4 FILLER_0_6_336 ();
 sg13g2_fill_2 FILLER_0_6_345 ();
 sg13g2_fill_1 FILLER_0_6_347 ();
 sg13g2_fill_2 FILLER_0_6_352 ();
 sg13g2_fill_2 FILLER_0_6_359 ();
 sg13g2_fill_8 FILLER_0_6_387 ();
 sg13g2_fill_8 FILLER_0_6_395 ();
 sg13g2_fill_8 FILLER_0_6_403 ();
 sg13g2_fill_1 FILLER_0_6_411 ();
 sg13g2_fill_2 FILLER_0_6_417 ();
 sg13g2_fill_1 FILLER_0_6_419 ();
 sg13g2_fill_8 FILLER_0_6_424 ();
 sg13g2_fill_8 FILLER_0_6_432 ();
 sg13g2_fill_4 FILLER_0_6_440 ();
 sg13g2_fill_1 FILLER_0_6_444 ();
 sg13g2_fill_2 FILLER_0_6_450 ();
 sg13g2_fill_8 FILLER_0_6_478 ();
 sg13g2_fill_8 FILLER_0_6_486 ();
 sg13g2_fill_8 FILLER_0_6_494 ();
 sg13g2_fill_8 FILLER_0_6_502 ();
 sg13g2_fill_2 FILLER_0_6_536 ();
 sg13g2_fill_2 FILLER_0_6_542 ();
 sg13g2_fill_2 FILLER_0_6_548 ();
 sg13g2_fill_1 FILLER_0_6_550 ();
 sg13g2_fill_8 FILLER_0_6_577 ();
 sg13g2_fill_8 FILLER_0_6_585 ();
 sg13g2_fill_4 FILLER_0_6_593 ();
 sg13g2_fill_2 FILLER_0_6_597 ();
 sg13g2_fill_1 FILLER_0_6_599 ();
 sg13g2_fill_2 FILLER_0_6_604 ();
 sg13g2_fill_8 FILLER_0_6_611 ();
 sg13g2_fill_8 FILLER_0_6_619 ();
 sg13g2_fill_8 FILLER_0_6_627 ();
 sg13g2_fill_8 FILLER_0_6_635 ();
 sg13g2_fill_8 FILLER_0_6_643 ();
 sg13g2_fill_8 FILLER_0_6_651 ();
 sg13g2_fill_8 FILLER_0_6_659 ();
 sg13g2_fill_4 FILLER_0_6_667 ();
 sg13g2_fill_2 FILLER_0_6_676 ();
 sg13g2_fill_2 FILLER_0_6_683 ();
 sg13g2_fill_2 FILLER_0_6_690 ();
 sg13g2_fill_8 FILLER_0_6_696 ();
 sg13g2_fill_8 FILLER_0_6_704 ();
 sg13g2_fill_8 FILLER_0_6_712 ();
 sg13g2_fill_4 FILLER_0_6_720 ();
 sg13g2_fill_2 FILLER_0_6_724 ();
 sg13g2_fill_2 FILLER_0_6_729 ();
 sg13g2_fill_4 FILLER_0_6_757 ();
 sg13g2_fill_2 FILLER_0_6_761 ();
 sg13g2_fill_1 FILLER_0_6_763 ();
 sg13g2_fill_8 FILLER_0_6_768 ();
 sg13g2_fill_1 FILLER_0_6_776 ();
 sg13g2_fill_2 FILLER_0_6_782 ();
 sg13g2_fill_2 FILLER_0_6_810 ();
 sg13g2_fill_8 FILLER_0_6_838 ();
 sg13g2_fill_4 FILLER_0_6_846 ();
 sg13g2_fill_2 FILLER_0_6_850 ();
 sg13g2_fill_1 FILLER_0_6_852 ();
 sg13g2_fill_2 FILLER_0_6_856 ();
 sg13g2_fill_8 FILLER_0_6_884 ();
 sg13g2_fill_8 FILLER_0_6_892 ();
 sg13g2_fill_8 FILLER_0_6_900 ();
 sg13g2_fill_2 FILLER_0_6_908 ();
 sg13g2_fill_8 FILLER_0_6_936 ();
 sg13g2_fill_8 FILLER_0_6_944 ();
 sg13g2_fill_8 FILLER_0_6_952 ();
 sg13g2_fill_8 FILLER_0_6_960 ();
 sg13g2_fill_4 FILLER_0_6_968 ();
 sg13g2_fill_2 FILLER_0_6_977 ();
 sg13g2_fill_8 FILLER_0_6_983 ();
 sg13g2_fill_8 FILLER_0_6_991 ();
 sg13g2_fill_4 FILLER_0_6_999 ();
 sg13g2_fill_1 FILLER_0_6_1003 ();
 sg13g2_fill_8 FILLER_0_6_1009 ();
 sg13g2_fill_8 FILLER_0_6_1017 ();
 sg13g2_fill_8 FILLER_0_6_1025 ();
 sg13g2_fill_8 FILLER_0_6_1033 ();
 sg13g2_fill_8 FILLER_0_6_1041 ();
 sg13g2_fill_1 FILLER_0_6_1049 ();
 sg13g2_fill_2 FILLER_0_6_1055 ();
 sg13g2_fill_4 FILLER_0_6_1083 ();
 sg13g2_fill_2 FILLER_0_6_1087 ();
 sg13g2_fill_1 FILLER_0_6_1089 ();
 sg13g2_fill_8 FILLER_0_6_1093 ();
 sg13g2_fill_4 FILLER_0_6_1101 ();
 sg13g2_fill_2 FILLER_0_6_1105 ();
 sg13g2_fill_1 FILLER_0_6_1107 ();
 sg13g2_fill_8 FILLER_0_6_1112 ();
 sg13g2_fill_8 FILLER_0_6_1120 ();
 sg13g2_fill_8 FILLER_0_6_1128 ();
 sg13g2_fill_8 FILLER_0_6_1136 ();
 sg13g2_fill_8 FILLER_0_6_1144 ();
 sg13g2_fill_8 FILLER_0_6_1152 ();
 sg13g2_fill_8 FILLER_0_6_1160 ();
 sg13g2_fill_8 FILLER_0_6_1168 ();
 sg13g2_fill_2 FILLER_0_6_1176 ();
 sg13g2_fill_1 FILLER_0_6_1178 ();
 sg13g2_fill_2 FILLER_0_6_1200 ();
 sg13g2_fill_8 FILLER_0_6_1228 ();
 sg13g2_fill_8 FILLER_0_6_1236 ();
 sg13g2_fill_8 FILLER_0_6_1244 ();
 sg13g2_fill_8 FILLER_0_6_1252 ();
 sg13g2_fill_8 FILLER_0_6_1260 ();
 sg13g2_fill_8 FILLER_0_6_1268 ();
 sg13g2_fill_8 FILLER_0_6_1276 ();
 sg13g2_fill_8 FILLER_0_6_1284 ();
 sg13g2_fill_4 FILLER_0_6_1292 ();
 sg13g2_fill_1 FILLER_0_6_1296 ();
 sg13g2_fill_8 FILLER_0_7_0 ();
 sg13g2_fill_8 FILLER_0_7_8 ();
 sg13g2_fill_8 FILLER_0_7_16 ();
 sg13g2_fill_8 FILLER_0_7_24 ();
 sg13g2_fill_8 FILLER_0_7_32 ();
 sg13g2_fill_8 FILLER_0_7_40 ();
 sg13g2_fill_8 FILLER_0_7_48 ();
 sg13g2_fill_8 FILLER_0_7_56 ();
 sg13g2_fill_8 FILLER_0_7_64 ();
 sg13g2_fill_8 FILLER_0_7_72 ();
 sg13g2_fill_8 FILLER_0_7_80 ();
 sg13g2_fill_8 FILLER_0_7_88 ();
 sg13g2_fill_8 FILLER_0_7_96 ();
 sg13g2_fill_8 FILLER_0_7_104 ();
 sg13g2_fill_8 FILLER_0_7_112 ();
 sg13g2_fill_8 FILLER_0_7_120 ();
 sg13g2_fill_8 FILLER_0_7_128 ();
 sg13g2_fill_8 FILLER_0_7_136 ();
 sg13g2_fill_8 FILLER_0_7_144 ();
 sg13g2_fill_8 FILLER_0_7_152 ();
 sg13g2_fill_8 FILLER_0_7_160 ();
 sg13g2_fill_8 FILLER_0_7_168 ();
 sg13g2_fill_8 FILLER_0_7_176 ();
 sg13g2_fill_8 FILLER_0_7_184 ();
 sg13g2_fill_8 FILLER_0_7_192 ();
 sg13g2_fill_8 FILLER_0_7_200 ();
 sg13g2_fill_8 FILLER_0_7_208 ();
 sg13g2_fill_8 FILLER_0_7_216 ();
 sg13g2_fill_8 FILLER_0_7_224 ();
 sg13g2_fill_8 FILLER_0_7_232 ();
 sg13g2_fill_8 FILLER_0_7_240 ();
 sg13g2_fill_8 FILLER_0_7_248 ();
 sg13g2_fill_8 FILLER_0_7_256 ();
 sg13g2_fill_8 FILLER_0_7_264 ();
 sg13g2_fill_8 FILLER_0_7_272 ();
 sg13g2_fill_8 FILLER_0_7_280 ();
 sg13g2_fill_8 FILLER_0_7_288 ();
 sg13g2_fill_8 FILLER_0_7_296 ();
 sg13g2_fill_8 FILLER_0_7_304 ();
 sg13g2_fill_8 FILLER_0_7_312 ();
 sg13g2_fill_8 FILLER_0_7_320 ();
 sg13g2_fill_8 FILLER_0_7_328 ();
 sg13g2_fill_2 FILLER_0_7_336 ();
 sg13g2_fill_1 FILLER_0_7_338 ();
 sg13g2_fill_4 FILLER_0_7_365 ();
 sg13g2_fill_2 FILLER_0_7_369 ();
 sg13g2_fill_8 FILLER_0_7_397 ();
 sg13g2_fill_8 FILLER_0_7_405 ();
 sg13g2_fill_4 FILLER_0_7_439 ();
 sg13g2_fill_2 FILLER_0_7_443 ();
 sg13g2_fill_1 FILLER_0_7_445 ();
 sg13g2_fill_2 FILLER_0_7_467 ();
 sg13g2_fill_8 FILLER_0_7_473 ();
 sg13g2_fill_8 FILLER_0_7_481 ();
 sg13g2_fill_8 FILLER_0_7_489 ();
 sg13g2_fill_4 FILLER_0_7_497 ();
 sg13g2_fill_1 FILLER_0_7_501 ();
 sg13g2_fill_2 FILLER_0_7_507 ();
 sg13g2_fill_4 FILLER_0_7_513 ();
 sg13g2_fill_2 FILLER_0_7_517 ();
 sg13g2_fill_2 FILLER_0_7_545 ();
 sg13g2_fill_1 FILLER_0_7_547 ();
 sg13g2_fill_2 FILLER_0_7_569 ();
 sg13g2_fill_1 FILLER_0_7_571 ();
 sg13g2_fill_2 FILLER_0_7_577 ();
 sg13g2_fill_1 FILLER_0_7_579 ();
 sg13g2_fill_4 FILLER_0_7_606 ();
 sg13g2_fill_8 FILLER_0_7_636 ();
 sg13g2_fill_8 FILLER_0_7_644 ();
 sg13g2_fill_8 FILLER_0_7_652 ();
 sg13g2_fill_1 FILLER_0_7_660 ();
 sg13g2_fill_2 FILLER_0_7_666 ();
 sg13g2_fill_2 FILLER_0_7_694 ();
 sg13g2_fill_1 FILLER_0_7_696 ();
 sg13g2_fill_4 FILLER_0_7_702 ();
 sg13g2_fill_2 FILLER_0_7_711 ();
 sg13g2_fill_2 FILLER_0_7_717 ();
 sg13g2_fill_8 FILLER_0_7_745 ();
 sg13g2_fill_8 FILLER_0_7_753 ();
 sg13g2_fill_2 FILLER_0_7_761 ();
 sg13g2_fill_4 FILLER_0_7_768 ();
 sg13g2_fill_2 FILLER_0_7_772 ();
 sg13g2_fill_1 FILLER_0_7_774 ();
 sg13g2_fill_2 FILLER_0_7_801 ();
 sg13g2_fill_2 FILLER_0_7_808 ();
 sg13g2_fill_2 FILLER_0_7_814 ();
 sg13g2_fill_2 FILLER_0_7_837 ();
 sg13g2_fill_8 FILLER_0_7_844 ();
 sg13g2_fill_8 FILLER_0_7_852 ();
 sg13g2_fill_2 FILLER_0_7_865 ();
 sg13g2_fill_1 FILLER_0_7_867 ();
 sg13g2_fill_4 FILLER_0_7_872 ();
 sg13g2_fill_2 FILLER_0_7_876 ();
 sg13g2_fill_1 FILLER_0_7_878 ();
 sg13g2_fill_2 FILLER_0_7_884 ();
 sg13g2_fill_8 FILLER_0_7_890 ();
 sg13g2_fill_2 FILLER_0_7_898 ();
 sg13g2_fill_1 FILLER_0_7_900 ();
 sg13g2_fill_4 FILLER_0_7_927 ();
 sg13g2_fill_8 FILLER_0_7_935 ();
 sg13g2_fill_8 FILLER_0_7_943 ();
 sg13g2_fill_8 FILLER_0_7_951 ();
 sg13g2_fill_2 FILLER_0_7_963 ();
 sg13g2_fill_1 FILLER_0_7_965 ();
 sg13g2_fill_4 FILLER_0_7_992 ();
 sg13g2_fill_2 FILLER_0_7_1000 ();
 sg13g2_fill_1 FILLER_0_7_1002 ();
 sg13g2_fill_8 FILLER_0_7_1007 ();
 sg13g2_fill_8 FILLER_0_7_1015 ();
 sg13g2_fill_1 FILLER_0_7_1023 ();
 sg13g2_fill_8 FILLER_0_7_1045 ();
 sg13g2_fill_8 FILLER_0_7_1053 ();
 sg13g2_fill_8 FILLER_0_7_1065 ();
 sg13g2_fill_4 FILLER_0_7_1073 ();
 sg13g2_fill_2 FILLER_0_7_1077 ();
 sg13g2_fill_1 FILLER_0_7_1079 ();
 sg13g2_fill_8 FILLER_0_7_1084 ();
 sg13g2_fill_8 FILLER_0_7_1092 ();
 sg13g2_fill_4 FILLER_0_7_1100 ();
 sg13g2_fill_2 FILLER_0_7_1104 ();
 sg13g2_fill_1 FILLER_0_7_1106 ();
 sg13g2_fill_2 FILLER_0_7_1112 ();
 sg13g2_fill_8 FILLER_0_7_1140 ();
 sg13g2_fill_8 FILLER_0_7_1148 ();
 sg13g2_fill_8 FILLER_0_7_1156 ();
 sg13g2_fill_8 FILLER_0_7_1164 ();
 sg13g2_fill_2 FILLER_0_7_1172 ();
 sg13g2_fill_1 FILLER_0_7_1174 ();
 sg13g2_fill_2 FILLER_0_7_1201 ();
 sg13g2_fill_4 FILLER_0_7_1207 ();
 sg13g2_fill_2 FILLER_0_7_1211 ();
 sg13g2_fill_1 FILLER_0_7_1213 ();
 sg13g2_fill_4 FILLER_0_7_1219 ();
 sg13g2_fill_2 FILLER_0_7_1223 ();
 sg13g2_fill_8 FILLER_0_7_1229 ();
 sg13g2_fill_8 FILLER_0_7_1237 ();
 sg13g2_fill_8 FILLER_0_7_1245 ();
 sg13g2_fill_8 FILLER_0_7_1253 ();
 sg13g2_fill_8 FILLER_0_7_1261 ();
 sg13g2_fill_8 FILLER_0_7_1269 ();
 sg13g2_fill_8 FILLER_0_7_1277 ();
 sg13g2_fill_8 FILLER_0_7_1285 ();
 sg13g2_fill_4 FILLER_0_7_1293 ();
 sg13g2_fill_8 FILLER_0_8_0 ();
 sg13g2_fill_8 FILLER_0_8_8 ();
 sg13g2_fill_8 FILLER_0_8_16 ();
 sg13g2_fill_8 FILLER_0_8_24 ();
 sg13g2_fill_8 FILLER_0_8_32 ();
 sg13g2_fill_8 FILLER_0_8_40 ();
 sg13g2_fill_8 FILLER_0_8_48 ();
 sg13g2_fill_8 FILLER_0_8_56 ();
 sg13g2_fill_8 FILLER_0_8_64 ();
 sg13g2_fill_8 FILLER_0_8_72 ();
 sg13g2_fill_8 FILLER_0_8_80 ();
 sg13g2_fill_8 FILLER_0_8_88 ();
 sg13g2_fill_8 FILLER_0_8_96 ();
 sg13g2_fill_8 FILLER_0_8_104 ();
 sg13g2_fill_8 FILLER_0_8_112 ();
 sg13g2_fill_8 FILLER_0_8_120 ();
 sg13g2_fill_8 FILLER_0_8_128 ();
 sg13g2_fill_8 FILLER_0_8_136 ();
 sg13g2_fill_8 FILLER_0_8_144 ();
 sg13g2_fill_8 FILLER_0_8_152 ();
 sg13g2_fill_8 FILLER_0_8_160 ();
 sg13g2_fill_8 FILLER_0_8_168 ();
 sg13g2_fill_8 FILLER_0_8_176 ();
 sg13g2_fill_8 FILLER_0_8_184 ();
 sg13g2_fill_8 FILLER_0_8_192 ();
 sg13g2_fill_8 FILLER_0_8_200 ();
 sg13g2_fill_8 FILLER_0_8_208 ();
 sg13g2_fill_8 FILLER_0_8_216 ();
 sg13g2_fill_8 FILLER_0_8_224 ();
 sg13g2_fill_8 FILLER_0_8_232 ();
 sg13g2_fill_8 FILLER_0_8_240 ();
 sg13g2_fill_8 FILLER_0_8_248 ();
 sg13g2_fill_8 FILLER_0_8_256 ();
 sg13g2_fill_8 FILLER_0_8_264 ();
 sg13g2_fill_8 FILLER_0_8_272 ();
 sg13g2_fill_8 FILLER_0_8_280 ();
 sg13g2_fill_8 FILLER_0_8_288 ();
 sg13g2_fill_8 FILLER_0_8_296 ();
 sg13g2_fill_8 FILLER_0_8_304 ();
 sg13g2_fill_8 FILLER_0_8_312 ();
 sg13g2_fill_4 FILLER_0_8_320 ();
 sg13g2_fill_1 FILLER_0_8_324 ();
 sg13g2_fill_8 FILLER_0_8_330 ();
 sg13g2_fill_4 FILLER_0_8_338 ();
 sg13g2_fill_1 FILLER_0_8_342 ();
 sg13g2_fill_8 FILLER_0_8_347 ();
 sg13g2_fill_4 FILLER_0_8_355 ();
 sg13g2_fill_2 FILLER_0_8_359 ();
 sg13g2_fill_2 FILLER_0_8_371 ();
 sg13g2_fill_4 FILLER_0_8_378 ();
 sg13g2_fill_1 FILLER_0_8_382 ();
 sg13g2_fill_8 FILLER_0_8_404 ();
 sg13g2_fill_4 FILLER_0_8_412 ();
 sg13g2_fill_1 FILLER_0_8_416 ();
 sg13g2_fill_2 FILLER_0_8_422 ();
 sg13g2_fill_4 FILLER_0_8_428 ();
 sg13g2_fill_2 FILLER_0_8_458 ();
 sg13g2_fill_8 FILLER_0_8_464 ();
 sg13g2_fill_8 FILLER_0_8_472 ();
 sg13g2_fill_4 FILLER_0_8_480 ();
 sg13g2_fill_2 FILLER_0_8_484 ();
 sg13g2_fill_1 FILLER_0_8_486 ();
 sg13g2_fill_8 FILLER_0_8_491 ();
 sg13g2_fill_8 FILLER_0_8_499 ();
 sg13g2_fill_8 FILLER_0_8_507 ();
 sg13g2_fill_4 FILLER_0_8_515 ();
 sg13g2_fill_2 FILLER_0_8_519 ();
 sg13g2_fill_2 FILLER_0_8_526 ();
 sg13g2_fill_2 FILLER_0_8_532 ();
 sg13g2_fill_8 FILLER_0_8_555 ();
 sg13g2_fill_8 FILLER_0_8_563 ();
 sg13g2_fill_4 FILLER_0_8_571 ();
 sg13g2_fill_2 FILLER_0_8_580 ();
 sg13g2_fill_2 FILLER_0_8_608 ();
 sg13g2_fill_1 FILLER_0_8_610 ();
 sg13g2_fill_4 FILLER_0_8_615 ();
 sg13g2_fill_1 FILLER_0_8_619 ();
 sg13g2_fill_2 FILLER_0_8_641 ();
 sg13g2_fill_2 FILLER_0_8_648 ();
 sg13g2_fill_1 FILLER_0_8_650 ();
 sg13g2_fill_2 FILLER_0_8_656 ();
 sg13g2_fill_8 FILLER_0_8_662 ();
 sg13g2_fill_2 FILLER_0_8_670 ();
 sg13g2_fill_1 FILLER_0_8_672 ();
 sg13g2_fill_2 FILLER_0_8_677 ();
 sg13g2_fill_2 FILLER_0_8_705 ();
 sg13g2_fill_8 FILLER_0_8_713 ();
 sg13g2_fill_8 FILLER_0_8_721 ();
 sg13g2_fill_4 FILLER_0_8_729 ();
 sg13g2_fill_2 FILLER_0_8_738 ();
 sg13g2_fill_2 FILLER_0_8_744 ();
 sg13g2_fill_8 FILLER_0_8_756 ();
 sg13g2_fill_8 FILLER_0_8_764 ();
 sg13g2_fill_8 FILLER_0_8_772 ();
 sg13g2_fill_8 FILLER_0_8_780 ();
 sg13g2_fill_1 FILLER_0_8_788 ();
 sg13g2_fill_2 FILLER_0_8_793 ();
 sg13g2_fill_8 FILLER_0_8_800 ();
 sg13g2_fill_1 FILLER_0_8_808 ();
 sg13g2_fill_4 FILLER_0_8_830 ();
 sg13g2_fill_1 FILLER_0_8_834 ();
 sg13g2_fill_2 FILLER_0_8_840 ();
 sg13g2_fill_4 FILLER_0_8_846 ();
 sg13g2_fill_2 FILLER_0_8_850 ();
 sg13g2_fill_4 FILLER_0_8_857 ();
 sg13g2_fill_2 FILLER_0_8_866 ();
 sg13g2_fill_4 FILLER_0_8_894 ();
 sg13g2_fill_2 FILLER_0_8_903 ();
 sg13g2_fill_2 FILLER_0_8_909 ();
 sg13g2_fill_1 FILLER_0_8_911 ();
 sg13g2_fill_4 FILLER_0_8_917 ();
 sg13g2_fill_1 FILLER_0_8_921 ();
 sg13g2_fill_2 FILLER_0_8_926 ();
 sg13g2_fill_8 FILLER_0_8_933 ();
 sg13g2_fill_8 FILLER_0_8_941 ();
 sg13g2_fill_8 FILLER_0_8_949 ();
 sg13g2_fill_2 FILLER_0_8_957 ();
 sg13g2_fill_8 FILLER_0_8_964 ();
 sg13g2_fill_4 FILLER_0_8_972 ();
 sg13g2_fill_2 FILLER_0_8_997 ();
 sg13g2_fill_2 FILLER_0_8_1004 ();
 sg13g2_fill_8 FILLER_0_8_1032 ();
 sg13g2_fill_2 FILLER_0_8_1040 ();
 sg13g2_fill_1 FILLER_0_8_1042 ();
 sg13g2_fill_8 FILLER_0_8_1048 ();
 sg13g2_fill_8 FILLER_0_8_1056 ();
 sg13g2_fill_8 FILLER_0_8_1064 ();
 sg13g2_fill_8 FILLER_0_8_1072 ();
 sg13g2_fill_1 FILLER_0_8_1080 ();
 sg13g2_fill_2 FILLER_0_8_1086 ();
 sg13g2_fill_4 FILLER_0_8_1092 ();
 sg13g2_fill_1 FILLER_0_8_1096 ();
 sg13g2_fill_2 FILLER_0_8_1102 ();
 sg13g2_fill_4 FILLER_0_8_1130 ();
 sg13g2_fill_2 FILLER_0_8_1155 ();
 sg13g2_fill_8 FILLER_0_8_1162 ();
 sg13g2_fill_4 FILLER_0_8_1175 ();
 sg13g2_fill_4 FILLER_0_8_1183 ();
 sg13g2_fill_1 FILLER_0_8_1187 ();
 sg13g2_fill_4 FILLER_0_8_1193 ();
 sg13g2_fill_1 FILLER_0_8_1197 ();
 sg13g2_fill_8 FILLER_0_8_1219 ();
 sg13g2_fill_8 FILLER_0_8_1227 ();
 sg13g2_fill_8 FILLER_0_8_1235 ();
 sg13g2_fill_8 FILLER_0_8_1243 ();
 sg13g2_fill_8 FILLER_0_8_1251 ();
 sg13g2_fill_8 FILLER_0_8_1259 ();
 sg13g2_fill_8 FILLER_0_8_1267 ();
 sg13g2_fill_8 FILLER_0_8_1275 ();
 sg13g2_fill_8 FILLER_0_8_1283 ();
 sg13g2_fill_4 FILLER_0_8_1291 ();
 sg13g2_fill_2 FILLER_0_8_1295 ();
 sg13g2_fill_8 FILLER_0_9_0 ();
 sg13g2_fill_8 FILLER_0_9_8 ();
 sg13g2_fill_8 FILLER_0_9_16 ();
 sg13g2_fill_8 FILLER_0_9_24 ();
 sg13g2_fill_8 FILLER_0_9_32 ();
 sg13g2_fill_8 FILLER_0_9_40 ();
 sg13g2_fill_8 FILLER_0_9_48 ();
 sg13g2_fill_8 FILLER_0_9_56 ();
 sg13g2_fill_8 FILLER_0_9_64 ();
 sg13g2_fill_8 FILLER_0_9_72 ();
 sg13g2_fill_8 FILLER_0_9_80 ();
 sg13g2_fill_8 FILLER_0_9_88 ();
 sg13g2_fill_8 FILLER_0_9_96 ();
 sg13g2_fill_8 FILLER_0_9_104 ();
 sg13g2_fill_8 FILLER_0_9_112 ();
 sg13g2_fill_8 FILLER_0_9_120 ();
 sg13g2_fill_8 FILLER_0_9_128 ();
 sg13g2_fill_8 FILLER_0_9_136 ();
 sg13g2_fill_8 FILLER_0_9_144 ();
 sg13g2_fill_8 FILLER_0_9_152 ();
 sg13g2_fill_8 FILLER_0_9_160 ();
 sg13g2_fill_8 FILLER_0_9_168 ();
 sg13g2_fill_8 FILLER_0_9_176 ();
 sg13g2_fill_8 FILLER_0_9_184 ();
 sg13g2_fill_8 FILLER_0_9_192 ();
 sg13g2_fill_8 FILLER_0_9_200 ();
 sg13g2_fill_8 FILLER_0_9_208 ();
 sg13g2_fill_8 FILLER_0_9_216 ();
 sg13g2_fill_8 FILLER_0_9_224 ();
 sg13g2_fill_8 FILLER_0_9_232 ();
 sg13g2_fill_8 FILLER_0_9_240 ();
 sg13g2_fill_8 FILLER_0_9_248 ();
 sg13g2_fill_8 FILLER_0_9_256 ();
 sg13g2_fill_8 FILLER_0_9_264 ();
 sg13g2_fill_8 FILLER_0_9_272 ();
 sg13g2_fill_8 FILLER_0_9_280 ();
 sg13g2_fill_8 FILLER_0_9_288 ();
 sg13g2_fill_8 FILLER_0_9_296 ();
 sg13g2_fill_8 FILLER_0_9_304 ();
 sg13g2_fill_8 FILLER_0_9_312 ();
 sg13g2_fill_1 FILLER_0_9_320 ();
 sg13g2_fill_8 FILLER_0_9_347 ();
 sg13g2_fill_8 FILLER_0_9_355 ();
 sg13g2_fill_8 FILLER_0_9_363 ();
 sg13g2_fill_8 FILLER_0_9_371 ();
 sg13g2_fill_2 FILLER_0_9_383 ();
 sg13g2_fill_8 FILLER_0_9_390 ();
 sg13g2_fill_8 FILLER_0_9_398 ();
 sg13g2_fill_8 FILLER_0_9_406 ();
 sg13g2_fill_8 FILLER_0_9_414 ();
 sg13g2_fill_8 FILLER_0_9_422 ();
 sg13g2_fill_8 FILLER_0_9_430 ();
 sg13g2_fill_4 FILLER_0_9_438 ();
 sg13g2_fill_8 FILLER_0_9_445 ();
 sg13g2_fill_8 FILLER_0_9_453 ();
 sg13g2_fill_8 FILLER_0_9_461 ();
 sg13g2_fill_8 FILLER_0_9_469 ();
 sg13g2_fill_8 FILLER_0_9_477 ();
 sg13g2_fill_4 FILLER_0_9_485 ();
 sg13g2_fill_2 FILLER_0_9_489 ();
 sg13g2_fill_2 FILLER_0_9_496 ();
 sg13g2_fill_8 FILLER_0_9_503 ();
 sg13g2_fill_8 FILLER_0_9_511 ();
 sg13g2_fill_8 FILLER_0_9_519 ();
 sg13g2_fill_8 FILLER_0_9_527 ();
 sg13g2_fill_8 FILLER_0_9_535 ();
 sg13g2_fill_8 FILLER_0_9_543 ();
 sg13g2_fill_2 FILLER_0_9_556 ();
 sg13g2_fill_8 FILLER_0_9_563 ();
 sg13g2_fill_8 FILLER_0_9_571 ();
 sg13g2_fill_8 FILLER_0_9_579 ();
 sg13g2_fill_2 FILLER_0_9_587 ();
 sg13g2_fill_8 FILLER_0_9_594 ();
 sg13g2_fill_2 FILLER_0_9_602 ();
 sg13g2_fill_4 FILLER_0_9_608 ();
 sg13g2_fill_1 FILLER_0_9_612 ();
 sg13g2_fill_8 FILLER_0_9_634 ();
 sg13g2_fill_8 FILLER_0_9_668 ();
 sg13g2_fill_4 FILLER_0_9_681 ();
 sg13g2_fill_2 FILLER_0_9_685 ();
 sg13g2_fill_8 FILLER_0_9_708 ();
 sg13g2_fill_8 FILLER_0_9_716 ();
 sg13g2_fill_8 FILLER_0_9_724 ();
 sg13g2_fill_8 FILLER_0_9_732 ();
 sg13g2_fill_8 FILLER_0_9_740 ();
 sg13g2_fill_8 FILLER_0_9_748 ();
 sg13g2_fill_8 FILLER_0_9_756 ();
 sg13g2_fill_8 FILLER_0_9_764 ();
 sg13g2_fill_8 FILLER_0_9_772 ();
 sg13g2_fill_4 FILLER_0_9_780 ();
 sg13g2_fill_2 FILLER_0_9_784 ();
 sg13g2_fill_2 FILLER_0_9_791 ();
 sg13g2_fill_2 FILLER_0_9_819 ();
 sg13g2_fill_8 FILLER_0_9_826 ();
 sg13g2_fill_8 FILLER_0_9_834 ();
 sg13g2_fill_2 FILLER_0_9_842 ();
 sg13g2_fill_2 FILLER_0_9_848 ();
 sg13g2_fill_8 FILLER_0_9_855 ();
 sg13g2_fill_8 FILLER_0_9_863 ();
 sg13g2_fill_4 FILLER_0_9_871 ();
 sg13g2_fill_2 FILLER_0_9_875 ();
 sg13g2_fill_8 FILLER_0_9_883 ();
 sg13g2_fill_8 FILLER_0_9_891 ();
 sg13g2_fill_1 FILLER_0_9_899 ();
 sg13g2_fill_8 FILLER_0_9_905 ();
 sg13g2_fill_1 FILLER_0_9_913 ();
 sg13g2_fill_8 FILLER_0_9_919 ();
 sg13g2_fill_2 FILLER_0_9_927 ();
 sg13g2_fill_1 FILLER_0_9_929 ();
 sg13g2_fill_8 FILLER_0_9_936 ();
 sg13g2_fill_8 FILLER_0_9_944 ();
 sg13g2_fill_4 FILLER_0_9_952 ();
 sg13g2_fill_8 FILLER_0_9_982 ();
 sg13g2_fill_8 FILLER_0_9_990 ();
 sg13g2_fill_2 FILLER_0_9_998 ();
 sg13g2_fill_2 FILLER_0_9_1008 ();
 sg13g2_fill_2 FILLER_0_9_1015 ();
 sg13g2_fill_8 FILLER_0_9_1021 ();
 sg13g2_fill_8 FILLER_0_9_1029 ();
 sg13g2_fill_8 FILLER_0_9_1037 ();
 sg13g2_fill_2 FILLER_0_9_1045 ();
 sg13g2_fill_1 FILLER_0_9_1047 ();
 sg13g2_fill_2 FILLER_0_9_1053 ();
 sg13g2_fill_8 FILLER_0_9_1059 ();
 sg13g2_fill_8 FILLER_0_9_1067 ();
 sg13g2_fill_8 FILLER_0_9_1075 ();
 sg13g2_fill_8 FILLER_0_9_1083 ();
 sg13g2_fill_8 FILLER_0_9_1091 ();
 sg13g2_fill_8 FILLER_0_9_1099 ();
 sg13g2_fill_2 FILLER_0_9_1107 ();
 sg13g2_fill_1 FILLER_0_9_1109 ();
 sg13g2_fill_2 FILLER_0_9_1114 ();
 sg13g2_fill_4 FILLER_0_9_1126 ();
 sg13g2_fill_2 FILLER_0_9_1130 ();
 sg13g2_fill_1 FILLER_0_9_1132 ();
 sg13g2_fill_2 FILLER_0_9_1159 ();
 sg13g2_fill_8 FILLER_0_9_1165 ();
 sg13g2_fill_8 FILLER_0_9_1173 ();
 sg13g2_fill_2 FILLER_0_9_1181 ();
 sg13g2_fill_1 FILLER_0_9_1183 ();
 sg13g2_fill_8 FILLER_0_9_1188 ();
 sg13g2_fill_8 FILLER_0_9_1196 ();
 sg13g2_fill_8 FILLER_0_9_1204 ();
 sg13g2_fill_8 FILLER_0_9_1212 ();
 sg13g2_fill_8 FILLER_0_9_1220 ();
 sg13g2_fill_8 FILLER_0_9_1228 ();
 sg13g2_fill_8 FILLER_0_9_1236 ();
 sg13g2_fill_8 FILLER_0_9_1244 ();
 sg13g2_fill_8 FILLER_0_9_1252 ();
 sg13g2_fill_8 FILLER_0_9_1260 ();
 sg13g2_fill_8 FILLER_0_9_1268 ();
 sg13g2_fill_8 FILLER_0_9_1276 ();
 sg13g2_fill_8 FILLER_0_9_1284 ();
 sg13g2_fill_4 FILLER_0_9_1292 ();
 sg13g2_fill_1 FILLER_0_9_1296 ();
 sg13g2_fill_8 FILLER_0_10_0 ();
 sg13g2_fill_8 FILLER_0_10_8 ();
 sg13g2_fill_8 FILLER_0_10_16 ();
 sg13g2_fill_8 FILLER_0_10_24 ();
 sg13g2_fill_8 FILLER_0_10_32 ();
 sg13g2_fill_8 FILLER_0_10_40 ();
 sg13g2_fill_8 FILLER_0_10_48 ();
 sg13g2_fill_8 FILLER_0_10_56 ();
 sg13g2_fill_8 FILLER_0_10_64 ();
 sg13g2_fill_8 FILLER_0_10_72 ();
 sg13g2_fill_8 FILLER_0_10_80 ();
 sg13g2_fill_8 FILLER_0_10_88 ();
 sg13g2_fill_8 FILLER_0_10_96 ();
 sg13g2_fill_8 FILLER_0_10_104 ();
 sg13g2_fill_8 FILLER_0_10_112 ();
 sg13g2_fill_8 FILLER_0_10_120 ();
 sg13g2_fill_8 FILLER_0_10_128 ();
 sg13g2_fill_8 FILLER_0_10_136 ();
 sg13g2_fill_8 FILLER_0_10_144 ();
 sg13g2_fill_8 FILLER_0_10_152 ();
 sg13g2_fill_8 FILLER_0_10_160 ();
 sg13g2_fill_8 FILLER_0_10_168 ();
 sg13g2_fill_8 FILLER_0_10_176 ();
 sg13g2_fill_8 FILLER_0_10_184 ();
 sg13g2_fill_8 FILLER_0_10_192 ();
 sg13g2_fill_8 FILLER_0_10_200 ();
 sg13g2_fill_8 FILLER_0_10_208 ();
 sg13g2_fill_8 FILLER_0_10_216 ();
 sg13g2_fill_8 FILLER_0_10_224 ();
 sg13g2_fill_8 FILLER_0_10_232 ();
 sg13g2_fill_8 FILLER_0_10_240 ();
 sg13g2_fill_8 FILLER_0_10_248 ();
 sg13g2_fill_8 FILLER_0_10_256 ();
 sg13g2_fill_8 FILLER_0_10_264 ();
 sg13g2_fill_8 FILLER_0_10_272 ();
 sg13g2_fill_8 FILLER_0_10_280 ();
 sg13g2_fill_8 FILLER_0_10_288 ();
 sg13g2_fill_8 FILLER_0_10_296 ();
 sg13g2_fill_8 FILLER_0_10_304 ();
 sg13g2_fill_8 FILLER_0_10_312 ();
 sg13g2_fill_8 FILLER_0_10_320 ();
 sg13g2_fill_8 FILLER_0_10_328 ();
 sg13g2_fill_2 FILLER_0_10_336 ();
 sg13g2_fill_2 FILLER_0_10_343 ();
 sg13g2_fill_2 FILLER_0_10_349 ();
 sg13g2_fill_2 FILLER_0_10_356 ();
 sg13g2_fill_4 FILLER_0_10_364 ();
 sg13g2_fill_1 FILLER_0_10_368 ();
 sg13g2_fill_2 FILLER_0_10_374 ();
 sg13g2_fill_8 FILLER_0_10_402 ();
 sg13g2_fill_8 FILLER_0_10_410 ();
 sg13g2_fill_8 FILLER_0_10_418 ();
 sg13g2_fill_8 FILLER_0_10_426 ();
 sg13g2_fill_8 FILLER_0_10_434 ();
 sg13g2_fill_4 FILLER_0_10_442 ();
 sg13g2_fill_2 FILLER_0_10_446 ();
 sg13g2_fill_2 FILLER_0_10_453 ();
 sg13g2_fill_8 FILLER_0_10_476 ();
 sg13g2_fill_1 FILLER_0_10_484 ();
 sg13g2_fill_8 FILLER_0_10_511 ();
 sg13g2_fill_8 FILLER_0_10_519 ();
 sg13g2_fill_8 FILLER_0_10_527 ();
 sg13g2_fill_8 FILLER_0_10_535 ();
 sg13g2_fill_8 FILLER_0_10_543 ();
 sg13g2_fill_8 FILLER_0_10_551 ();
 sg13g2_fill_4 FILLER_0_10_559 ();
 sg13g2_fill_2 FILLER_0_10_563 ();
 sg13g2_fill_8 FILLER_0_10_571 ();
 sg13g2_fill_8 FILLER_0_10_579 ();
 sg13g2_fill_8 FILLER_0_10_587 ();
 sg13g2_fill_8 FILLER_0_10_595 ();
 sg13g2_fill_8 FILLER_0_10_603 ();
 sg13g2_fill_8 FILLER_0_10_611 ();
 sg13g2_fill_8 FILLER_0_10_619 ();
 sg13g2_fill_8 FILLER_0_10_637 ();
 sg13g2_fill_2 FILLER_0_10_650 ();
 sg13g2_fill_8 FILLER_0_10_678 ();
 sg13g2_fill_2 FILLER_0_10_686 ();
 sg13g2_fill_1 FILLER_0_10_688 ();
 sg13g2_fill_8 FILLER_0_10_694 ();
 sg13g2_fill_2 FILLER_0_10_702 ();
 sg13g2_fill_2 FILLER_0_10_709 ();
 sg13g2_fill_8 FILLER_0_10_719 ();
 sg13g2_fill_8 FILLER_0_10_727 ();
 sg13g2_fill_8 FILLER_0_10_735 ();
 sg13g2_fill_8 FILLER_0_10_743 ();
 sg13g2_fill_8 FILLER_0_10_751 ();
 sg13g2_fill_8 FILLER_0_10_759 ();
 sg13g2_fill_8 FILLER_0_10_767 ();
 sg13g2_fill_4 FILLER_0_10_775 ();
 sg13g2_fill_1 FILLER_0_10_779 ();
 sg13g2_fill_8 FILLER_0_10_785 ();
 sg13g2_fill_8 FILLER_0_10_793 ();
 sg13g2_fill_4 FILLER_0_10_801 ();
 sg13g2_fill_8 FILLER_0_10_810 ();
 sg13g2_fill_1 FILLER_0_10_818 ();
 sg13g2_fill_8 FILLER_0_10_823 ();
 sg13g2_fill_1 FILLER_0_10_831 ();
 sg13g2_fill_8 FILLER_0_10_837 ();
 sg13g2_fill_8 FILLER_0_10_845 ();
 sg13g2_fill_8 FILLER_0_10_853 ();
 sg13g2_fill_8 FILLER_0_10_861 ();
 sg13g2_fill_8 FILLER_0_10_869 ();
 sg13g2_fill_8 FILLER_0_10_877 ();
 sg13g2_fill_8 FILLER_0_10_885 ();
 sg13g2_fill_8 FILLER_0_10_893 ();
 sg13g2_fill_8 FILLER_0_10_901 ();
 sg13g2_fill_4 FILLER_0_10_909 ();
 sg13g2_fill_1 FILLER_0_10_913 ();
 sg13g2_fill_8 FILLER_0_10_917 ();
 sg13g2_fill_8 FILLER_0_10_925 ();
 sg13g2_fill_8 FILLER_0_10_933 ();
 sg13g2_fill_8 FILLER_0_10_941 ();
 sg13g2_fill_8 FILLER_0_10_949 ();
 sg13g2_fill_8 FILLER_0_10_957 ();
 sg13g2_fill_8 FILLER_0_10_965 ();
 sg13g2_fill_8 FILLER_0_10_973 ();
 sg13g2_fill_2 FILLER_0_10_981 ();
 sg13g2_fill_1 FILLER_0_10_983 ();
 sg13g2_fill_8 FILLER_0_10_988 ();
 sg13g2_fill_4 FILLER_0_10_996 ();
 sg13g2_fill_2 FILLER_0_10_1000 ();
 sg13g2_fill_1 FILLER_0_10_1002 ();
 sg13g2_fill_2 FILLER_0_10_1008 ();
 sg13g2_fill_4 FILLER_0_10_1036 ();
 sg13g2_fill_2 FILLER_0_10_1040 ();
 sg13g2_fill_1 FILLER_0_10_1042 ();
 sg13g2_fill_8 FILLER_0_10_1069 ();
 sg13g2_fill_8 FILLER_0_10_1077 ();
 sg13g2_fill_8 FILLER_0_10_1085 ();
 sg13g2_fill_8 FILLER_0_10_1093 ();
 sg13g2_fill_8 FILLER_0_10_1101 ();
 sg13g2_fill_8 FILLER_0_10_1109 ();
 sg13g2_fill_8 FILLER_0_10_1117 ();
 sg13g2_fill_4 FILLER_0_10_1125 ();
 sg13g2_fill_2 FILLER_0_10_1129 ();
 sg13g2_fill_8 FILLER_0_10_1157 ();
 sg13g2_fill_8 FILLER_0_10_1165 ();
 sg13g2_fill_8 FILLER_0_10_1173 ();
 sg13g2_fill_2 FILLER_0_10_1181 ();
 sg13g2_fill_1 FILLER_0_10_1183 ();
 sg13g2_fill_2 FILLER_0_10_1189 ();
 sg13g2_fill_8 FILLER_0_10_1217 ();
 sg13g2_fill_8 FILLER_0_10_1225 ();
 sg13g2_fill_8 FILLER_0_10_1233 ();
 sg13g2_fill_8 FILLER_0_10_1241 ();
 sg13g2_fill_8 FILLER_0_10_1249 ();
 sg13g2_fill_8 FILLER_0_10_1257 ();
 sg13g2_fill_8 FILLER_0_10_1265 ();
 sg13g2_fill_8 FILLER_0_10_1273 ();
 sg13g2_fill_8 FILLER_0_10_1281 ();
 sg13g2_fill_8 FILLER_0_10_1289 ();
 sg13g2_fill_8 FILLER_0_11_0 ();
 sg13g2_fill_8 FILLER_0_11_8 ();
 sg13g2_fill_8 FILLER_0_11_16 ();
 sg13g2_fill_8 FILLER_0_11_24 ();
 sg13g2_fill_8 FILLER_0_11_32 ();
 sg13g2_fill_8 FILLER_0_11_40 ();
 sg13g2_fill_8 FILLER_0_11_48 ();
 sg13g2_fill_8 FILLER_0_11_56 ();
 sg13g2_fill_8 FILLER_0_11_64 ();
 sg13g2_fill_8 FILLER_0_11_72 ();
 sg13g2_fill_8 FILLER_0_11_80 ();
 sg13g2_fill_8 FILLER_0_11_88 ();
 sg13g2_fill_8 FILLER_0_11_96 ();
 sg13g2_fill_8 FILLER_0_11_104 ();
 sg13g2_fill_8 FILLER_0_11_112 ();
 sg13g2_fill_8 FILLER_0_11_120 ();
 sg13g2_fill_8 FILLER_0_11_128 ();
 sg13g2_fill_8 FILLER_0_11_136 ();
 sg13g2_fill_8 FILLER_0_11_144 ();
 sg13g2_fill_8 FILLER_0_11_152 ();
 sg13g2_fill_8 FILLER_0_11_160 ();
 sg13g2_fill_8 FILLER_0_11_168 ();
 sg13g2_fill_8 FILLER_0_11_176 ();
 sg13g2_fill_8 FILLER_0_11_184 ();
 sg13g2_fill_8 FILLER_0_11_192 ();
 sg13g2_fill_8 FILLER_0_11_200 ();
 sg13g2_fill_8 FILLER_0_11_208 ();
 sg13g2_fill_8 FILLER_0_11_216 ();
 sg13g2_fill_8 FILLER_0_11_224 ();
 sg13g2_fill_8 FILLER_0_11_232 ();
 sg13g2_fill_8 FILLER_0_11_240 ();
 sg13g2_fill_8 FILLER_0_11_248 ();
 sg13g2_fill_8 FILLER_0_11_256 ();
 sg13g2_fill_8 FILLER_0_11_264 ();
 sg13g2_fill_8 FILLER_0_11_272 ();
 sg13g2_fill_8 FILLER_0_11_280 ();
 sg13g2_fill_2 FILLER_0_11_288 ();
 sg13g2_fill_4 FILLER_0_11_316 ();
 sg13g2_fill_4 FILLER_0_11_324 ();
 sg13g2_fill_2 FILLER_0_11_328 ();
 sg13g2_fill_2 FILLER_0_11_356 ();
 sg13g2_fill_4 FILLER_0_11_364 ();
 sg13g2_fill_1 FILLER_0_11_368 ();
 sg13g2_fill_4 FILLER_0_11_375 ();
 sg13g2_fill_2 FILLER_0_11_379 ();
 sg13g2_fill_8 FILLER_0_11_387 ();
 sg13g2_fill_1 FILLER_0_11_395 ();
 sg13g2_fill_8 FILLER_0_11_400 ();
 sg13g2_fill_2 FILLER_0_11_413 ();
 sg13g2_fill_1 FILLER_0_11_415 ();
 sg13g2_fill_2 FILLER_0_11_420 ();
 sg13g2_fill_8 FILLER_0_11_432 ();
 sg13g2_fill_4 FILLER_0_11_440 ();
 sg13g2_fill_2 FILLER_0_11_444 ();
 sg13g2_fill_8 FILLER_0_11_451 ();
 sg13g2_fill_2 FILLER_0_11_459 ();
 sg13g2_fill_4 FILLER_0_11_471 ();
 sg13g2_fill_2 FILLER_0_11_475 ();
 sg13g2_fill_1 FILLER_0_11_477 ();
 sg13g2_fill_2 FILLER_0_11_483 ();
 sg13g2_fill_8 FILLER_0_11_489 ();
 sg13g2_fill_8 FILLER_0_11_497 ();
 sg13g2_fill_8 FILLER_0_11_510 ();
 sg13g2_fill_8 FILLER_0_11_518 ();
 sg13g2_fill_4 FILLER_0_11_526 ();
 sg13g2_fill_8 FILLER_0_11_556 ();
 sg13g2_fill_8 FILLER_0_11_564 ();
 sg13g2_fill_8 FILLER_0_11_572 ();
 sg13g2_fill_2 FILLER_0_11_580 ();
 sg13g2_fill_1 FILLER_0_11_582 ();
 sg13g2_fill_2 FILLER_0_11_588 ();
 sg13g2_fill_8 FILLER_0_11_598 ();
 sg13g2_fill_8 FILLER_0_11_606 ();
 sg13g2_fill_8 FILLER_0_11_614 ();
 sg13g2_fill_8 FILLER_0_11_622 ();
 sg13g2_fill_8 FILLER_0_11_630 ();
 sg13g2_fill_8 FILLER_0_11_638 ();
 sg13g2_fill_8 FILLER_0_11_646 ();
 sg13g2_fill_1 FILLER_0_11_654 ();
 sg13g2_fill_2 FILLER_0_11_660 ();
 sg13g2_fill_4 FILLER_0_11_666 ();
 sg13g2_fill_1 FILLER_0_11_670 ();
 sg13g2_fill_2 FILLER_0_11_676 ();
 sg13g2_fill_8 FILLER_0_11_684 ();
 sg13g2_fill_8 FILLER_0_11_692 ();
 sg13g2_fill_8 FILLER_0_11_700 ();
 sg13g2_fill_8 FILLER_0_11_708 ();
 sg13g2_fill_8 FILLER_0_11_716 ();
 sg13g2_fill_2 FILLER_0_11_724 ();
 sg13g2_fill_1 FILLER_0_11_726 ();
 sg13g2_fill_4 FILLER_0_11_732 ();
 sg13g2_fill_2 FILLER_0_11_740 ();
 sg13g2_fill_4 FILLER_0_11_746 ();
 sg13g2_fill_2 FILLER_0_11_750 ();
 sg13g2_fill_2 FILLER_0_11_773 ();
 sg13g2_fill_8 FILLER_0_11_801 ();
 sg13g2_fill_8 FILLER_0_11_809 ();
 sg13g2_fill_8 FILLER_0_11_817 ();
 sg13g2_fill_4 FILLER_0_11_825 ();
 sg13g2_fill_2 FILLER_0_11_829 ();
 sg13g2_fill_1 FILLER_0_11_831 ();
 sg13g2_fill_4 FILLER_0_11_836 ();
 sg13g2_fill_2 FILLER_0_11_840 ();
 sg13g2_fill_1 FILLER_0_11_842 ();
 sg13g2_fill_2 FILLER_0_11_848 ();
 sg13g2_fill_4 FILLER_0_11_854 ();
 sg13g2_fill_2 FILLER_0_11_858 ();
 sg13g2_fill_2 FILLER_0_11_864 ();
 sg13g2_fill_2 FILLER_0_11_871 ();
 sg13g2_fill_8 FILLER_0_11_878 ();
 sg13g2_fill_8 FILLER_0_11_886 ();
 sg13g2_fill_8 FILLER_0_11_894 ();
 sg13g2_fill_8 FILLER_0_11_902 ();
 sg13g2_fill_4 FILLER_0_11_910 ();
 sg13g2_fill_2 FILLER_0_11_914 ();
 sg13g2_fill_4 FILLER_0_11_921 ();
 sg13g2_fill_2 FILLER_0_11_925 ();
 sg13g2_fill_1 FILLER_0_11_927 ();
 sg13g2_fill_8 FILLER_0_11_934 ();
 sg13g2_fill_8 FILLER_0_11_942 ();
 sg13g2_fill_8 FILLER_0_11_950 ();
 sg13g2_fill_8 FILLER_0_11_958 ();
 sg13g2_fill_1 FILLER_0_11_966 ();
 sg13g2_fill_8 FILLER_0_11_993 ();
 sg13g2_fill_4 FILLER_0_11_1001 ();
 sg13g2_fill_1 FILLER_0_11_1005 ();
 sg13g2_fill_8 FILLER_0_11_1010 ();
 sg13g2_fill_1 FILLER_0_11_1018 ();
 sg13g2_fill_8 FILLER_0_11_1029 ();
 sg13g2_fill_8 FILLER_0_11_1037 ();
 sg13g2_fill_8 FILLER_0_11_1045 ();
 sg13g2_fill_4 FILLER_0_11_1053 ();
 sg13g2_fill_4 FILLER_0_11_1062 ();
 sg13g2_fill_2 FILLER_0_11_1066 ();
 sg13g2_fill_1 FILLER_0_11_1068 ();
 sg13g2_fill_2 FILLER_0_11_1073 ();
 sg13g2_fill_4 FILLER_0_11_1085 ();
 sg13g2_fill_8 FILLER_0_11_1110 ();
 sg13g2_fill_8 FILLER_0_11_1118 ();
 sg13g2_fill_2 FILLER_0_11_1126 ();
 sg13g2_fill_2 FILLER_0_11_1133 ();
 sg13g2_fill_1 FILLER_0_11_1135 ();
 sg13g2_fill_2 FILLER_0_11_1140 ();
 sg13g2_fill_8 FILLER_0_11_1152 ();
 sg13g2_fill_8 FILLER_0_11_1160 ();
 sg13g2_fill_8 FILLER_0_11_1168 ();
 sg13g2_fill_8 FILLER_0_11_1176 ();
 sg13g2_fill_8 FILLER_0_11_1184 ();
 sg13g2_fill_8 FILLER_0_11_1192 ();
 sg13g2_fill_8 FILLER_0_11_1200 ();
 sg13g2_fill_8 FILLER_0_11_1208 ();
 sg13g2_fill_8 FILLER_0_11_1216 ();
 sg13g2_fill_8 FILLER_0_11_1224 ();
 sg13g2_fill_8 FILLER_0_11_1232 ();
 sg13g2_fill_8 FILLER_0_11_1240 ();
 sg13g2_fill_8 FILLER_0_11_1248 ();
 sg13g2_fill_8 FILLER_0_11_1256 ();
 sg13g2_fill_8 FILLER_0_11_1264 ();
 sg13g2_fill_8 FILLER_0_11_1272 ();
 sg13g2_fill_8 FILLER_0_11_1280 ();
 sg13g2_fill_8 FILLER_0_11_1288 ();
 sg13g2_fill_1 FILLER_0_11_1296 ();
 sg13g2_fill_8 FILLER_0_12_0 ();
 sg13g2_fill_8 FILLER_0_12_8 ();
 sg13g2_fill_8 FILLER_0_12_16 ();
 sg13g2_fill_8 FILLER_0_12_24 ();
 sg13g2_fill_8 FILLER_0_12_32 ();
 sg13g2_fill_8 FILLER_0_12_40 ();
 sg13g2_fill_8 FILLER_0_12_48 ();
 sg13g2_fill_8 FILLER_0_12_56 ();
 sg13g2_fill_8 FILLER_0_12_64 ();
 sg13g2_fill_8 FILLER_0_12_72 ();
 sg13g2_fill_8 FILLER_0_12_80 ();
 sg13g2_fill_8 FILLER_0_12_88 ();
 sg13g2_fill_8 FILLER_0_12_96 ();
 sg13g2_fill_8 FILLER_0_12_104 ();
 sg13g2_fill_8 FILLER_0_12_112 ();
 sg13g2_fill_8 FILLER_0_12_120 ();
 sg13g2_fill_8 FILLER_0_12_128 ();
 sg13g2_fill_8 FILLER_0_12_136 ();
 sg13g2_fill_8 FILLER_0_12_144 ();
 sg13g2_fill_8 FILLER_0_12_152 ();
 sg13g2_fill_8 FILLER_0_12_160 ();
 sg13g2_fill_8 FILLER_0_12_168 ();
 sg13g2_fill_8 FILLER_0_12_176 ();
 sg13g2_fill_8 FILLER_0_12_184 ();
 sg13g2_fill_8 FILLER_0_12_192 ();
 sg13g2_fill_8 FILLER_0_12_200 ();
 sg13g2_fill_8 FILLER_0_12_208 ();
 sg13g2_fill_8 FILLER_0_12_216 ();
 sg13g2_fill_8 FILLER_0_12_224 ();
 sg13g2_fill_8 FILLER_0_12_232 ();
 sg13g2_fill_8 FILLER_0_12_240 ();
 sg13g2_fill_8 FILLER_0_12_248 ();
 sg13g2_fill_8 FILLER_0_12_256 ();
 sg13g2_fill_8 FILLER_0_12_264 ();
 sg13g2_fill_8 FILLER_0_12_272 ();
 sg13g2_fill_8 FILLER_0_12_280 ();
 sg13g2_fill_8 FILLER_0_12_288 ();
 sg13g2_fill_4 FILLER_0_12_296 ();
 sg13g2_fill_2 FILLER_0_12_300 ();
 sg13g2_fill_2 FILLER_0_12_328 ();
 sg13g2_fill_8 FILLER_0_12_351 ();
 sg13g2_fill_8 FILLER_0_12_359 ();
 sg13g2_fill_8 FILLER_0_12_367 ();
 sg13g2_fill_8 FILLER_0_12_375 ();
 sg13g2_fill_8 FILLER_0_12_383 ();
 sg13g2_fill_1 FILLER_0_12_391 ();
 sg13g2_fill_8 FILLER_0_12_397 ();
 sg13g2_fill_8 FILLER_0_12_405 ();
 sg13g2_fill_4 FILLER_0_12_439 ();
 sg13g2_fill_4 FILLER_0_12_469 ();
 sg13g2_fill_1 FILLER_0_12_473 ();
 sg13g2_fill_8 FILLER_0_12_478 ();
 sg13g2_fill_8 FILLER_0_12_486 ();
 sg13g2_fill_2 FILLER_0_12_494 ();
 sg13g2_fill_1 FILLER_0_12_496 ();
 sg13g2_fill_4 FILLER_0_12_502 ();
 sg13g2_fill_2 FILLER_0_12_506 ();
 sg13g2_fill_1 FILLER_0_12_508 ();
 sg13g2_fill_8 FILLER_0_12_514 ();
 sg13g2_fill_8 FILLER_0_12_522 ();
 sg13g2_fill_1 FILLER_0_12_530 ();
 sg13g2_fill_4 FILLER_0_12_557 ();
 sg13g2_fill_1 FILLER_0_12_561 ();
 sg13g2_fill_2 FILLER_0_12_566 ();
 sg13g2_fill_4 FILLER_0_12_594 ();
 sg13g2_fill_8 FILLER_0_12_619 ();
 sg13g2_fill_8 FILLER_0_12_627 ();
 sg13g2_fill_8 FILLER_0_12_635 ();
 sg13g2_fill_8 FILLER_0_12_643 ();
 sg13g2_fill_8 FILLER_0_12_651 ();
 sg13g2_fill_8 FILLER_0_12_659 ();
 sg13g2_fill_8 FILLER_0_12_667 ();
 sg13g2_fill_8 FILLER_0_12_680 ();
 sg13g2_fill_8 FILLER_0_12_688 ();
 sg13g2_fill_8 FILLER_0_12_696 ();
 sg13g2_fill_8 FILLER_0_12_704 ();
 sg13g2_fill_8 FILLER_0_12_712 ();
 sg13g2_fill_4 FILLER_0_12_720 ();
 sg13g2_fill_1 FILLER_0_12_724 ();
 sg13g2_fill_2 FILLER_0_12_751 ();
 sg13g2_fill_4 FILLER_0_12_763 ();
 sg13g2_fill_1 FILLER_0_12_767 ();
 sg13g2_fill_2 FILLER_0_12_773 ();
 sg13g2_fill_2 FILLER_0_12_785 ();
 sg13g2_fill_8 FILLER_0_12_791 ();
 sg13g2_fill_8 FILLER_0_12_799 ();
 sg13g2_fill_4 FILLER_0_12_807 ();
 sg13g2_fill_1 FILLER_0_12_811 ();
 sg13g2_fill_2 FILLER_0_12_838 ();
 sg13g2_fill_2 FILLER_0_12_866 ();
 sg13g2_fill_2 FILLER_0_12_894 ();
 sg13g2_fill_1 FILLER_0_12_896 ();
 sg13g2_fill_2 FILLER_0_12_904 ();
 sg13g2_fill_1 FILLER_0_12_906 ();
 sg13g2_fill_4 FILLER_0_12_911 ();
 sg13g2_fill_8 FILLER_0_12_921 ();
 sg13g2_fill_1 FILLER_0_12_929 ();
 sg13g2_fill_4 FILLER_0_12_940 ();
 sg13g2_fill_2 FILLER_0_12_954 ();
 sg13g2_fill_1 FILLER_0_12_956 ();
 sg13g2_fill_2 FILLER_0_12_983 ();
 sg13g2_fill_8 FILLER_0_12_990 ();
 sg13g2_fill_8 FILLER_0_12_998 ();
 sg13g2_fill_8 FILLER_0_12_1006 ();
 sg13g2_fill_8 FILLER_0_12_1014 ();
 sg13g2_fill_8 FILLER_0_12_1022 ();
 sg13g2_fill_4 FILLER_0_12_1030 ();
 sg13g2_fill_8 FILLER_0_12_1039 ();
 sg13g2_fill_8 FILLER_0_12_1047 ();
 sg13g2_fill_8 FILLER_0_12_1055 ();
 sg13g2_fill_4 FILLER_0_12_1063 ();
 sg13g2_fill_2 FILLER_0_12_1067 ();
 sg13g2_fill_2 FILLER_0_12_1074 ();
 sg13g2_fill_2 FILLER_0_12_1102 ();
 sg13g2_fill_2 FILLER_0_12_1109 ();
 sg13g2_fill_1 FILLER_0_12_1111 ();
 sg13g2_fill_4 FILLER_0_12_1117 ();
 sg13g2_fill_8 FILLER_0_12_1126 ();
 sg13g2_fill_1 FILLER_0_12_1134 ();
 sg13g2_fill_8 FILLER_0_12_1139 ();
 sg13g2_fill_8 FILLER_0_12_1147 ();
 sg13g2_fill_8 FILLER_0_12_1155 ();
 sg13g2_fill_8 FILLER_0_12_1163 ();
 sg13g2_fill_8 FILLER_0_12_1171 ();
 sg13g2_fill_8 FILLER_0_12_1179 ();
 sg13g2_fill_8 FILLER_0_12_1187 ();
 sg13g2_fill_4 FILLER_0_12_1195 ();
 sg13g2_fill_2 FILLER_0_12_1204 ();
 sg13g2_fill_8 FILLER_0_12_1211 ();
 sg13g2_fill_8 FILLER_0_12_1219 ();
 sg13g2_fill_8 FILLER_0_12_1227 ();
 sg13g2_fill_8 FILLER_0_12_1235 ();
 sg13g2_fill_8 FILLER_0_12_1243 ();
 sg13g2_fill_8 FILLER_0_12_1251 ();
 sg13g2_fill_8 FILLER_0_12_1259 ();
 sg13g2_fill_8 FILLER_0_12_1267 ();
 sg13g2_fill_8 FILLER_0_12_1275 ();
 sg13g2_fill_8 FILLER_0_12_1283 ();
 sg13g2_fill_4 FILLER_0_12_1291 ();
 sg13g2_fill_2 FILLER_0_12_1295 ();
 sg13g2_fill_8 FILLER_0_13_0 ();
 sg13g2_fill_8 FILLER_0_13_8 ();
 sg13g2_fill_8 FILLER_0_13_16 ();
 sg13g2_fill_8 FILLER_0_13_24 ();
 sg13g2_fill_8 FILLER_0_13_32 ();
 sg13g2_fill_8 FILLER_0_13_40 ();
 sg13g2_fill_8 FILLER_0_13_48 ();
 sg13g2_fill_8 FILLER_0_13_56 ();
 sg13g2_fill_8 FILLER_0_13_64 ();
 sg13g2_fill_8 FILLER_0_13_72 ();
 sg13g2_fill_8 FILLER_0_13_80 ();
 sg13g2_fill_8 FILLER_0_13_88 ();
 sg13g2_fill_8 FILLER_0_13_96 ();
 sg13g2_fill_8 FILLER_0_13_104 ();
 sg13g2_fill_8 FILLER_0_13_112 ();
 sg13g2_fill_8 FILLER_0_13_120 ();
 sg13g2_fill_8 FILLER_0_13_128 ();
 sg13g2_fill_8 FILLER_0_13_136 ();
 sg13g2_fill_8 FILLER_0_13_144 ();
 sg13g2_fill_8 FILLER_0_13_152 ();
 sg13g2_fill_8 FILLER_0_13_160 ();
 sg13g2_fill_8 FILLER_0_13_168 ();
 sg13g2_fill_8 FILLER_0_13_176 ();
 sg13g2_fill_8 FILLER_0_13_184 ();
 sg13g2_fill_8 FILLER_0_13_192 ();
 sg13g2_fill_8 FILLER_0_13_200 ();
 sg13g2_fill_8 FILLER_0_13_208 ();
 sg13g2_fill_8 FILLER_0_13_216 ();
 sg13g2_fill_8 FILLER_0_13_224 ();
 sg13g2_fill_8 FILLER_0_13_232 ();
 sg13g2_fill_8 FILLER_0_13_240 ();
 sg13g2_fill_8 FILLER_0_13_248 ();
 sg13g2_fill_8 FILLER_0_13_256 ();
 sg13g2_fill_8 FILLER_0_13_264 ();
 sg13g2_fill_8 FILLER_0_13_272 ();
 sg13g2_fill_8 FILLER_0_13_280 ();
 sg13g2_fill_8 FILLER_0_13_288 ();
 sg13g2_fill_4 FILLER_0_13_296 ();
 sg13g2_fill_1 FILLER_0_13_300 ();
 sg13g2_fill_2 FILLER_0_13_305 ();
 sg13g2_fill_8 FILLER_0_13_312 ();
 sg13g2_fill_1 FILLER_0_13_320 ();
 sg13g2_fill_2 FILLER_0_13_326 ();
 sg13g2_fill_8 FILLER_0_13_333 ();
 sg13g2_fill_8 FILLER_0_13_341 ();
 sg13g2_fill_4 FILLER_0_13_349 ();
 sg13g2_fill_2 FILLER_0_13_357 ();
 sg13g2_fill_2 FILLER_0_13_364 ();
 sg13g2_fill_1 FILLER_0_13_366 ();
 sg13g2_fill_2 FILLER_0_13_372 ();
 sg13g2_fill_4 FILLER_0_13_379 ();
 sg13g2_fill_2 FILLER_0_13_383 ();
 sg13g2_fill_4 FILLER_0_13_390 ();
 sg13g2_fill_2 FILLER_0_13_394 ();
 sg13g2_fill_8 FILLER_0_13_400 ();
 sg13g2_fill_8 FILLER_0_13_408 ();
 sg13g2_fill_8 FILLER_0_13_416 ();
 sg13g2_fill_1 FILLER_0_13_424 ();
 sg13g2_fill_8 FILLER_0_13_433 ();
 sg13g2_fill_8 FILLER_0_13_441 ();
 sg13g2_fill_2 FILLER_0_13_449 ();
 sg13g2_fill_2 FILLER_0_13_455 ();
 sg13g2_fill_2 FILLER_0_13_483 ();
 sg13g2_fill_4 FILLER_0_13_490 ();
 sg13g2_fill_2 FILLER_0_13_494 ();
 sg13g2_fill_1 FILLER_0_13_496 ();
 sg13g2_fill_4 FILLER_0_13_502 ();
 sg13g2_fill_8 FILLER_0_13_513 ();
 sg13g2_fill_4 FILLER_0_13_521 ();
 sg13g2_fill_2 FILLER_0_13_525 ();
 sg13g2_fill_2 FILLER_0_13_532 ();
 sg13g2_fill_4 FILLER_0_13_538 ();
 sg13g2_fill_2 FILLER_0_13_542 ();
 sg13g2_fill_1 FILLER_0_13_544 ();
 sg13g2_fill_4 FILLER_0_13_555 ();
 sg13g2_fill_2 FILLER_0_13_559 ();
 sg13g2_fill_8 FILLER_0_13_566 ();
 sg13g2_fill_1 FILLER_0_13_574 ();
 sg13g2_fill_2 FILLER_0_13_601 ();
 sg13g2_fill_2 FILLER_0_13_608 ();
 sg13g2_fill_2 FILLER_0_13_616 ();
 sg13g2_fill_1 FILLER_0_13_618 ();
 sg13g2_fill_8 FILLER_0_13_623 ();
 sg13g2_fill_8 FILLER_0_13_631 ();
 sg13g2_fill_8 FILLER_0_13_639 ();
 sg13g2_fill_4 FILLER_0_13_647 ();
 sg13g2_fill_8 FILLER_0_13_677 ();
 sg13g2_fill_4 FILLER_0_13_685 ();
 sg13g2_fill_2 FILLER_0_13_689 ();
 sg13g2_fill_8 FILLER_0_13_696 ();
 sg13g2_fill_2 FILLER_0_13_704 ();
 sg13g2_fill_8 FILLER_0_13_710 ();
 sg13g2_fill_8 FILLER_0_13_718 ();
 sg13g2_fill_1 FILLER_0_13_726 ();
 sg13g2_fill_8 FILLER_0_13_753 ();
 sg13g2_fill_8 FILLER_0_13_761 ();
 sg13g2_fill_8 FILLER_0_13_769 ();
 sg13g2_fill_1 FILLER_0_13_777 ();
 sg13g2_fill_8 FILLER_0_13_783 ();
 sg13g2_fill_8 FILLER_0_13_791 ();
 sg13g2_fill_4 FILLER_0_13_799 ();
 sg13g2_fill_2 FILLER_0_13_803 ();
 sg13g2_fill_2 FILLER_0_13_831 ();
 sg13g2_fill_2 FILLER_0_13_854 ();
 sg13g2_fill_8 FILLER_0_13_861 ();
 sg13g2_fill_8 FILLER_0_13_869 ();
 sg13g2_fill_8 FILLER_0_13_877 ();
 sg13g2_fill_2 FILLER_0_13_885 ();
 sg13g2_fill_1 FILLER_0_13_887 ();
 sg13g2_fill_4 FILLER_0_13_891 ();
 sg13g2_fill_2 FILLER_0_13_895 ();
 sg13g2_fill_1 FILLER_0_13_897 ();
 sg13g2_fill_2 FILLER_0_13_924 ();
 sg13g2_fill_2 FILLER_0_13_952 ();
 sg13g2_fill_2 FILLER_0_13_959 ();
 sg13g2_fill_1 FILLER_0_13_961 ();
 sg13g2_fill_2 FILLER_0_13_967 ();
 sg13g2_fill_4 FILLER_0_13_973 ();
 sg13g2_fill_1 FILLER_0_13_977 ();
 sg13g2_fill_8 FILLER_0_13_999 ();
 sg13g2_fill_8 FILLER_0_13_1007 ();
 sg13g2_fill_8 FILLER_0_13_1015 ();
 sg13g2_fill_8 FILLER_0_13_1023 ();
 sg13g2_fill_8 FILLER_0_13_1031 ();
 sg13g2_fill_8 FILLER_0_13_1039 ();
 sg13g2_fill_4 FILLER_0_13_1047 ();
 sg13g2_fill_1 FILLER_0_13_1051 ();
 sg13g2_fill_2 FILLER_0_13_1057 ();
 sg13g2_fill_2 FILLER_0_13_1064 ();
 sg13g2_fill_2 FILLER_0_13_1071 ();
 sg13g2_fill_4 FILLER_0_13_1077 ();
 sg13g2_fill_2 FILLER_0_13_1081 ();
 sg13g2_fill_1 FILLER_0_13_1083 ();
 sg13g2_fill_2 FILLER_0_13_1089 ();
 sg13g2_fill_2 FILLER_0_13_1101 ();
 sg13g2_fill_8 FILLER_0_13_1107 ();
 sg13g2_fill_4 FILLER_0_13_1115 ();
 sg13g2_fill_2 FILLER_0_13_1119 ();
 sg13g2_fill_1 FILLER_0_13_1121 ();
 sg13g2_fill_8 FILLER_0_13_1148 ();
 sg13g2_fill_4 FILLER_0_13_1156 ();
 sg13g2_fill_2 FILLER_0_13_1160 ();
 sg13g2_fill_1 FILLER_0_13_1162 ();
 sg13g2_fill_8 FILLER_0_13_1168 ();
 sg13g2_fill_8 FILLER_0_13_1176 ();
 sg13g2_fill_8 FILLER_0_13_1184 ();
 sg13g2_fill_8 FILLER_0_13_1192 ();
 sg13g2_fill_2 FILLER_0_13_1200 ();
 sg13g2_fill_8 FILLER_0_13_1206 ();
 sg13g2_fill_8 FILLER_0_13_1214 ();
 sg13g2_fill_8 FILLER_0_13_1222 ();
 sg13g2_fill_8 FILLER_0_13_1230 ();
 sg13g2_fill_8 FILLER_0_13_1238 ();
 sg13g2_fill_8 FILLER_0_13_1246 ();
 sg13g2_fill_8 FILLER_0_13_1254 ();
 sg13g2_fill_8 FILLER_0_13_1262 ();
 sg13g2_fill_8 FILLER_0_13_1270 ();
 sg13g2_fill_8 FILLER_0_13_1278 ();
 sg13g2_fill_8 FILLER_0_13_1286 ();
 sg13g2_fill_2 FILLER_0_13_1294 ();
 sg13g2_fill_1 FILLER_0_13_1296 ();
 sg13g2_fill_8 FILLER_0_14_0 ();
 sg13g2_fill_8 FILLER_0_14_8 ();
 sg13g2_fill_8 FILLER_0_14_16 ();
 sg13g2_fill_8 FILLER_0_14_24 ();
 sg13g2_fill_8 FILLER_0_14_32 ();
 sg13g2_fill_8 FILLER_0_14_40 ();
 sg13g2_fill_8 FILLER_0_14_48 ();
 sg13g2_fill_8 FILLER_0_14_56 ();
 sg13g2_fill_8 FILLER_0_14_64 ();
 sg13g2_fill_8 FILLER_0_14_72 ();
 sg13g2_fill_8 FILLER_0_14_80 ();
 sg13g2_fill_8 FILLER_0_14_88 ();
 sg13g2_fill_8 FILLER_0_14_96 ();
 sg13g2_fill_8 FILLER_0_14_104 ();
 sg13g2_fill_8 FILLER_0_14_112 ();
 sg13g2_fill_8 FILLER_0_14_120 ();
 sg13g2_fill_8 FILLER_0_14_128 ();
 sg13g2_fill_8 FILLER_0_14_136 ();
 sg13g2_fill_8 FILLER_0_14_144 ();
 sg13g2_fill_8 FILLER_0_14_152 ();
 sg13g2_fill_8 FILLER_0_14_160 ();
 sg13g2_fill_8 FILLER_0_14_168 ();
 sg13g2_fill_8 FILLER_0_14_176 ();
 sg13g2_fill_8 FILLER_0_14_184 ();
 sg13g2_fill_8 FILLER_0_14_192 ();
 sg13g2_fill_8 FILLER_0_14_200 ();
 sg13g2_fill_8 FILLER_0_14_208 ();
 sg13g2_fill_8 FILLER_0_14_216 ();
 sg13g2_fill_8 FILLER_0_14_224 ();
 sg13g2_fill_8 FILLER_0_14_232 ();
 sg13g2_fill_8 FILLER_0_14_240 ();
 sg13g2_fill_8 FILLER_0_14_248 ();
 sg13g2_fill_8 FILLER_0_14_256 ();
 sg13g2_fill_8 FILLER_0_14_264 ();
 sg13g2_fill_8 FILLER_0_14_272 ();
 sg13g2_fill_8 FILLER_0_14_280 ();
 sg13g2_fill_8 FILLER_0_14_288 ();
 sg13g2_fill_8 FILLER_0_14_296 ();
 sg13g2_fill_8 FILLER_0_14_304 ();
 sg13g2_fill_8 FILLER_0_14_312 ();
 sg13g2_fill_8 FILLER_0_14_320 ();
 sg13g2_fill_8 FILLER_0_14_328 ();
 sg13g2_fill_8 FILLER_0_14_336 ();
 sg13g2_fill_2 FILLER_0_14_348 ();
 sg13g2_fill_2 FILLER_0_14_376 ();
 sg13g2_fill_2 FILLER_0_14_383 ();
 sg13g2_fill_2 FILLER_0_14_390 ();
 sg13g2_fill_2 FILLER_0_14_397 ();
 sg13g2_fill_8 FILLER_0_14_403 ();
 sg13g2_fill_8 FILLER_0_14_411 ();
 sg13g2_fill_4 FILLER_0_14_419 ();
 sg13g2_fill_2 FILLER_0_14_423 ();
 sg13g2_fill_1 FILLER_0_14_425 ();
 sg13g2_fill_4 FILLER_0_14_431 ();
 sg13g2_fill_2 FILLER_0_14_435 ();
 sg13g2_fill_1 FILLER_0_14_437 ();
 sg13g2_fill_2 FILLER_0_14_445 ();
 sg13g2_fill_8 FILLER_0_14_455 ();
 sg13g2_fill_8 FILLER_0_14_463 ();
 sg13g2_fill_8 FILLER_0_14_471 ();
 sg13g2_fill_4 FILLER_0_14_479 ();
 sg13g2_fill_2 FILLER_0_14_483 ();
 sg13g2_fill_2 FILLER_0_14_490 ();
 sg13g2_fill_2 FILLER_0_14_498 ();
 sg13g2_fill_8 FILLER_0_14_505 ();
 sg13g2_fill_8 FILLER_0_14_513 ();
 sg13g2_fill_8 FILLER_0_14_521 ();
 sg13g2_fill_4 FILLER_0_14_529 ();
 sg13g2_fill_1 FILLER_0_14_533 ();
 sg13g2_fill_4 FILLER_0_14_539 ();
 sg13g2_fill_1 FILLER_0_14_543 ();
 sg13g2_fill_8 FILLER_0_14_548 ();
 sg13g2_fill_8 FILLER_0_14_561 ();
 sg13g2_fill_8 FILLER_0_14_569 ();
 sg13g2_fill_2 FILLER_0_14_577 ();
 sg13g2_fill_4 FILLER_0_14_584 ();
 sg13g2_fill_2 FILLER_0_14_588 ();
 sg13g2_fill_1 FILLER_0_14_590 ();
 sg13g2_fill_8 FILLER_0_14_595 ();
 sg13g2_fill_1 FILLER_0_14_603 ();
 sg13g2_fill_2 FILLER_0_14_610 ();
 sg13g2_fill_2 FILLER_0_14_617 ();
 sg13g2_fill_2 FILLER_0_14_624 ();
 sg13g2_fill_8 FILLER_0_14_652 ();
 sg13g2_fill_2 FILLER_0_14_660 ();
 sg13g2_fill_1 FILLER_0_14_662 ();
 sg13g2_fill_2 FILLER_0_14_668 ();
 sg13g2_fill_1 FILLER_0_14_670 ();
 sg13g2_fill_2 FILLER_0_14_676 ();
 sg13g2_fill_1 FILLER_0_14_678 ();
 sg13g2_fill_2 FILLER_0_14_689 ();
 sg13g2_fill_8 FILLER_0_14_717 ();
 sg13g2_fill_8 FILLER_0_14_725 ();
 sg13g2_fill_4 FILLER_0_14_733 ();
 sg13g2_fill_2 FILLER_0_14_737 ();
 sg13g2_fill_2 FILLER_0_14_744 ();
 sg13g2_fill_8 FILLER_0_14_751 ();
 sg13g2_fill_8 FILLER_0_14_759 ();
 sg13g2_fill_1 FILLER_0_14_767 ();
 sg13g2_fill_8 FILLER_0_14_776 ();
 sg13g2_fill_4 FILLER_0_14_784 ();
 sg13g2_fill_2 FILLER_0_14_788 ();
 sg13g2_fill_8 FILLER_0_14_795 ();
 sg13g2_fill_4 FILLER_0_14_803 ();
 sg13g2_fill_2 FILLER_0_14_807 ();
 sg13g2_fill_2 FILLER_0_14_814 ();
 sg13g2_fill_2 FILLER_0_14_820 ();
 sg13g2_fill_8 FILLER_0_14_827 ();
 sg13g2_fill_2 FILLER_0_14_835 ();
 sg13g2_fill_2 FILLER_0_14_842 ();
 sg13g2_fill_2 FILLER_0_14_865 ();
 sg13g2_fill_8 FILLER_0_14_872 ();
 sg13g2_fill_2 FILLER_0_14_880 ();
 sg13g2_fill_1 FILLER_0_14_882 ();
 sg13g2_fill_2 FILLER_0_14_888 ();
 sg13g2_fill_1 FILLER_0_14_890 ();
 sg13g2_fill_8 FILLER_0_14_896 ();
 sg13g2_fill_4 FILLER_0_14_909 ();
 sg13g2_fill_2 FILLER_0_14_913 ();
 sg13g2_fill_8 FILLER_0_14_920 ();
 sg13g2_fill_4 FILLER_0_14_928 ();
 sg13g2_fill_2 FILLER_0_14_937 ();
 sg13g2_fill_8 FILLER_0_14_943 ();
 sg13g2_fill_8 FILLER_0_14_951 ();
 sg13g2_fill_8 FILLER_0_14_959 ();
 sg13g2_fill_8 FILLER_0_14_967 ();
 sg13g2_fill_8 FILLER_0_14_975 ();
 sg13g2_fill_2 FILLER_0_14_983 ();
 sg13g2_fill_2 FILLER_0_14_1006 ();
 sg13g2_fill_2 FILLER_0_14_1016 ();
 sg13g2_fill_2 FILLER_0_14_1023 ();
 sg13g2_fill_2 FILLER_0_14_1051 ();
 sg13g2_fill_1 FILLER_0_14_1053 ();
 sg13g2_fill_2 FILLER_0_14_1060 ();
 sg13g2_fill_2 FILLER_0_14_1067 ();
 sg13g2_fill_4 FILLER_0_14_1074 ();
 sg13g2_fill_8 FILLER_0_14_1104 ();
 sg13g2_fill_8 FILLER_0_14_1112 ();
 sg13g2_fill_8 FILLER_0_14_1120 ();
 sg13g2_fill_8 FILLER_0_14_1128 ();
 sg13g2_fill_4 FILLER_0_14_1136 ();
 sg13g2_fill_2 FILLER_0_14_1140 ();
 sg13g2_fill_8 FILLER_0_14_1145 ();
 sg13g2_fill_8 FILLER_0_14_1153 ();
 sg13g2_fill_8 FILLER_0_14_1161 ();
 sg13g2_fill_8 FILLER_0_14_1169 ();
 sg13g2_fill_8 FILLER_0_14_1177 ();
 sg13g2_fill_8 FILLER_0_14_1185 ();
 sg13g2_fill_4 FILLER_0_14_1193 ();
 sg13g2_fill_1 FILLER_0_14_1197 ();
 sg13g2_fill_8 FILLER_0_14_1224 ();
 sg13g2_fill_8 FILLER_0_14_1232 ();
 sg13g2_fill_8 FILLER_0_14_1240 ();
 sg13g2_fill_8 FILLER_0_14_1248 ();
 sg13g2_fill_8 FILLER_0_14_1256 ();
 sg13g2_fill_8 FILLER_0_14_1264 ();
 sg13g2_fill_8 FILLER_0_14_1272 ();
 sg13g2_fill_8 FILLER_0_14_1280 ();
 sg13g2_fill_8 FILLER_0_14_1288 ();
 sg13g2_fill_1 FILLER_0_14_1296 ();
 sg13g2_fill_8 FILLER_0_15_0 ();
 sg13g2_fill_8 FILLER_0_15_8 ();
 sg13g2_fill_8 FILLER_0_15_16 ();
 sg13g2_fill_8 FILLER_0_15_24 ();
 sg13g2_fill_8 FILLER_0_15_32 ();
 sg13g2_fill_8 FILLER_0_15_40 ();
 sg13g2_fill_8 FILLER_0_15_48 ();
 sg13g2_fill_8 FILLER_0_15_56 ();
 sg13g2_fill_8 FILLER_0_15_64 ();
 sg13g2_fill_8 FILLER_0_15_72 ();
 sg13g2_fill_8 FILLER_0_15_80 ();
 sg13g2_fill_8 FILLER_0_15_88 ();
 sg13g2_fill_8 FILLER_0_15_96 ();
 sg13g2_fill_8 FILLER_0_15_104 ();
 sg13g2_fill_8 FILLER_0_15_112 ();
 sg13g2_fill_8 FILLER_0_15_120 ();
 sg13g2_fill_8 FILLER_0_15_128 ();
 sg13g2_fill_8 FILLER_0_15_136 ();
 sg13g2_fill_8 FILLER_0_15_144 ();
 sg13g2_fill_8 FILLER_0_15_152 ();
 sg13g2_fill_8 FILLER_0_15_160 ();
 sg13g2_fill_8 FILLER_0_15_168 ();
 sg13g2_fill_8 FILLER_0_15_176 ();
 sg13g2_fill_8 FILLER_0_15_184 ();
 sg13g2_fill_8 FILLER_0_15_192 ();
 sg13g2_fill_8 FILLER_0_15_200 ();
 sg13g2_fill_8 FILLER_0_15_208 ();
 sg13g2_fill_8 FILLER_0_15_216 ();
 sg13g2_fill_8 FILLER_0_15_224 ();
 sg13g2_fill_8 FILLER_0_15_232 ();
 sg13g2_fill_8 FILLER_0_15_240 ();
 sg13g2_fill_8 FILLER_0_15_248 ();
 sg13g2_fill_8 FILLER_0_15_256 ();
 sg13g2_fill_8 FILLER_0_15_264 ();
 sg13g2_fill_8 FILLER_0_15_272 ();
 sg13g2_fill_8 FILLER_0_15_280 ();
 sg13g2_fill_8 FILLER_0_15_288 ();
 sg13g2_fill_8 FILLER_0_15_296 ();
 sg13g2_fill_8 FILLER_0_15_304 ();
 sg13g2_fill_8 FILLER_0_15_312 ();
 sg13g2_fill_4 FILLER_0_15_320 ();
 sg13g2_fill_2 FILLER_0_15_324 ();
 sg13g2_fill_8 FILLER_0_15_331 ();
 sg13g2_fill_8 FILLER_0_15_339 ();
 sg13g2_fill_4 FILLER_0_15_352 ();
 sg13g2_fill_1 FILLER_0_15_356 ();
 sg13g2_fill_2 FILLER_0_15_362 ();
 sg13g2_fill_2 FILLER_0_15_390 ();
 sg13g2_fill_4 FILLER_0_15_396 ();
 sg13g2_fill_2 FILLER_0_15_400 ();
 sg13g2_fill_8 FILLER_0_15_410 ();
 sg13g2_fill_8 FILLER_0_15_418 ();
 sg13g2_fill_8 FILLER_0_15_426 ();
 sg13g2_fill_8 FILLER_0_15_437 ();
 sg13g2_fill_4 FILLER_0_15_445 ();
 sg13g2_fill_1 FILLER_0_15_449 ();
 sg13g2_fill_8 FILLER_0_15_454 ();
 sg13g2_fill_8 FILLER_0_15_462 ();
 sg13g2_fill_8 FILLER_0_15_470 ();
 sg13g2_fill_8 FILLER_0_15_478 ();
 sg13g2_fill_8 FILLER_0_15_486 ();
 sg13g2_fill_4 FILLER_0_15_494 ();
 sg13g2_fill_2 FILLER_0_15_498 ();
 sg13g2_fill_1 FILLER_0_15_500 ();
 sg13g2_fill_4 FILLER_0_15_506 ();
 sg13g2_fill_8 FILLER_0_15_514 ();
 sg13g2_fill_8 FILLER_0_15_527 ();
 sg13g2_fill_1 FILLER_0_15_535 ();
 sg13g2_fill_8 FILLER_0_15_557 ();
 sg13g2_fill_2 FILLER_0_15_565 ();
 sg13g2_fill_8 FILLER_0_15_572 ();
 sg13g2_fill_8 FILLER_0_15_580 ();
 sg13g2_fill_8 FILLER_0_15_588 ();
 sg13g2_fill_8 FILLER_0_15_596 ();
 sg13g2_fill_8 FILLER_0_15_604 ();
 sg13g2_fill_4 FILLER_0_15_612 ();
 sg13g2_fill_2 FILLER_0_15_616 ();
 sg13g2_fill_1 FILLER_0_15_618 ();
 sg13g2_fill_4 FILLER_0_15_627 ();
 sg13g2_fill_1 FILLER_0_15_631 ();
 sg13g2_fill_2 FILLER_0_15_637 ();
 sg13g2_fill_8 FILLER_0_15_644 ();
 sg13g2_fill_8 FILLER_0_15_652 ();
 sg13g2_fill_8 FILLER_0_15_660 ();
 sg13g2_fill_2 FILLER_0_15_668 ();
 sg13g2_fill_1 FILLER_0_15_670 ();
 sg13g2_fill_8 FILLER_0_15_675 ();
 sg13g2_fill_1 FILLER_0_15_683 ();
 sg13g2_fill_2 FILLER_0_15_689 ();
 sg13g2_fill_2 FILLER_0_15_695 ();
 sg13g2_fill_1 FILLER_0_15_697 ();
 sg13g2_fill_8 FILLER_0_15_703 ();
 sg13g2_fill_8 FILLER_0_15_711 ();
 sg13g2_fill_8 FILLER_0_15_719 ();
 sg13g2_fill_8 FILLER_0_15_727 ();
 sg13g2_fill_8 FILLER_0_15_735 ();
 sg13g2_fill_8 FILLER_0_15_743 ();
 sg13g2_fill_8 FILLER_0_15_751 ();
 sg13g2_fill_8 FILLER_0_15_759 ();
 sg13g2_fill_8 FILLER_0_15_767 ();
 sg13g2_fill_2 FILLER_0_15_775 ();
 sg13g2_fill_8 FILLER_0_15_782 ();
 sg13g2_fill_2 FILLER_0_15_790 ();
 sg13g2_fill_1 FILLER_0_15_792 ();
 sg13g2_fill_8 FILLER_0_15_798 ();
 sg13g2_fill_8 FILLER_0_15_806 ();
 sg13g2_fill_1 FILLER_0_15_814 ();
 sg13g2_fill_8 FILLER_0_15_820 ();
 sg13g2_fill_1 FILLER_0_15_828 ();
 sg13g2_fill_8 FILLER_0_15_833 ();
 sg13g2_fill_4 FILLER_0_15_841 ();
 sg13g2_fill_2 FILLER_0_15_845 ();
 sg13g2_fill_8 FILLER_0_15_852 ();
 sg13g2_fill_8 FILLER_0_15_860 ();
 sg13g2_fill_8 FILLER_0_15_868 ();
 sg13g2_fill_8 FILLER_0_15_876 ();
 sg13g2_fill_8 FILLER_0_15_884 ();
 sg13g2_fill_8 FILLER_0_15_892 ();
 sg13g2_fill_8 FILLER_0_15_900 ();
 sg13g2_fill_8 FILLER_0_15_908 ();
 sg13g2_fill_8 FILLER_0_15_920 ();
 sg13g2_fill_8 FILLER_0_15_928 ();
 sg13g2_fill_8 FILLER_0_15_936 ();
 sg13g2_fill_4 FILLER_0_15_949 ();
 sg13g2_fill_2 FILLER_0_15_953 ();
 sg13g2_fill_8 FILLER_0_15_960 ();
 sg13g2_fill_8 FILLER_0_15_968 ();
 sg13g2_fill_8 FILLER_0_15_976 ();
 sg13g2_fill_8 FILLER_0_15_984 ();
 sg13g2_fill_8 FILLER_0_15_992 ();
 sg13g2_fill_4 FILLER_0_15_1000 ();
 sg13g2_fill_2 FILLER_0_15_1004 ();
 sg13g2_fill_4 FILLER_0_15_1011 ();
 sg13g2_fill_1 FILLER_0_15_1015 ();
 sg13g2_fill_8 FILLER_0_15_1022 ();
 sg13g2_fill_8 FILLER_0_15_1030 ();
 sg13g2_fill_8 FILLER_0_15_1038 ();
 sg13g2_fill_4 FILLER_0_15_1046 ();
 sg13g2_fill_2 FILLER_0_15_1055 ();
 sg13g2_fill_8 FILLER_0_15_1064 ();
 sg13g2_fill_8 FILLER_0_15_1072 ();
 sg13g2_fill_2 FILLER_0_15_1080 ();
 sg13g2_fill_8 FILLER_0_15_1086 ();
 sg13g2_fill_8 FILLER_0_15_1094 ();
 sg13g2_fill_8 FILLER_0_15_1102 ();
 sg13g2_fill_8 FILLER_0_15_1110 ();
 sg13g2_fill_1 FILLER_0_15_1118 ();
 sg13g2_fill_2 FILLER_0_15_1124 ();
 sg13g2_fill_8 FILLER_0_15_1130 ();
 sg13g2_fill_8 FILLER_0_15_1138 ();
 sg13g2_fill_4 FILLER_0_15_1151 ();
 sg13g2_fill_2 FILLER_0_15_1155 ();
 sg13g2_fill_8 FILLER_0_15_1161 ();
 sg13g2_fill_8 FILLER_0_15_1169 ();
 sg13g2_fill_8 FILLER_0_15_1177 ();
 sg13g2_fill_2 FILLER_0_15_1185 ();
 sg13g2_fill_1 FILLER_0_15_1187 ();
 sg13g2_fill_2 FILLER_0_15_1193 ();
 sg13g2_fill_8 FILLER_0_15_1199 ();
 sg13g2_fill_4 FILLER_0_15_1207 ();
 sg13g2_fill_2 FILLER_0_15_1211 ();
 sg13g2_fill_8 FILLER_0_15_1234 ();
 sg13g2_fill_8 FILLER_0_15_1242 ();
 sg13g2_fill_8 FILLER_0_15_1250 ();
 sg13g2_fill_8 FILLER_0_15_1258 ();
 sg13g2_fill_8 FILLER_0_15_1266 ();
 sg13g2_fill_8 FILLER_0_15_1274 ();
 sg13g2_fill_8 FILLER_0_15_1282 ();
 sg13g2_fill_4 FILLER_0_15_1290 ();
 sg13g2_fill_2 FILLER_0_15_1294 ();
 sg13g2_fill_1 FILLER_0_15_1296 ();
 sg13g2_fill_8 FILLER_0_16_0 ();
 sg13g2_fill_8 FILLER_0_16_8 ();
 sg13g2_fill_8 FILLER_0_16_16 ();
 sg13g2_fill_8 FILLER_0_16_24 ();
 sg13g2_fill_8 FILLER_0_16_32 ();
 sg13g2_fill_8 FILLER_0_16_40 ();
 sg13g2_fill_8 FILLER_0_16_48 ();
 sg13g2_fill_8 FILLER_0_16_56 ();
 sg13g2_fill_8 FILLER_0_16_64 ();
 sg13g2_fill_8 FILLER_0_16_72 ();
 sg13g2_fill_8 FILLER_0_16_80 ();
 sg13g2_fill_8 FILLER_0_16_88 ();
 sg13g2_fill_8 FILLER_0_16_96 ();
 sg13g2_fill_8 FILLER_0_16_104 ();
 sg13g2_fill_8 FILLER_0_16_112 ();
 sg13g2_fill_8 FILLER_0_16_120 ();
 sg13g2_fill_8 FILLER_0_16_128 ();
 sg13g2_fill_8 FILLER_0_16_136 ();
 sg13g2_fill_8 FILLER_0_16_144 ();
 sg13g2_fill_8 FILLER_0_16_152 ();
 sg13g2_fill_8 FILLER_0_16_160 ();
 sg13g2_fill_8 FILLER_0_16_168 ();
 sg13g2_fill_8 FILLER_0_16_176 ();
 sg13g2_fill_8 FILLER_0_16_184 ();
 sg13g2_fill_8 FILLER_0_16_192 ();
 sg13g2_fill_8 FILLER_0_16_200 ();
 sg13g2_fill_8 FILLER_0_16_208 ();
 sg13g2_fill_8 FILLER_0_16_216 ();
 sg13g2_fill_8 FILLER_0_16_224 ();
 sg13g2_fill_8 FILLER_0_16_232 ();
 sg13g2_fill_8 FILLER_0_16_240 ();
 sg13g2_fill_8 FILLER_0_16_248 ();
 sg13g2_fill_8 FILLER_0_16_256 ();
 sg13g2_fill_8 FILLER_0_16_264 ();
 sg13g2_fill_8 FILLER_0_16_272 ();
 sg13g2_fill_8 FILLER_0_16_280 ();
 sg13g2_fill_8 FILLER_0_16_288 ();
 sg13g2_fill_4 FILLER_0_16_296 ();
 sg13g2_fill_1 FILLER_0_16_300 ();
 sg13g2_fill_8 FILLER_0_16_306 ();
 sg13g2_fill_1 FILLER_0_16_314 ();
 sg13g2_fill_8 FILLER_0_16_319 ();
 sg13g2_fill_4 FILLER_0_16_327 ();
 sg13g2_fill_2 FILLER_0_16_331 ();
 sg13g2_fill_1 FILLER_0_16_333 ();
 sg13g2_fill_8 FILLER_0_16_339 ();
 sg13g2_fill_4 FILLER_0_16_347 ();
 sg13g2_fill_2 FILLER_0_16_351 ();
 sg13g2_fill_2 FILLER_0_16_357 ();
 sg13g2_fill_2 FILLER_0_16_365 ();
 sg13g2_fill_2 FILLER_0_16_377 ();
 sg13g2_fill_4 FILLER_0_16_384 ();
 sg13g2_fill_2 FILLER_0_16_388 ();
 sg13g2_fill_1 FILLER_0_16_390 ();
 sg13g2_fill_8 FILLER_0_16_399 ();
 sg13g2_fill_8 FILLER_0_16_407 ();
 sg13g2_fill_8 FILLER_0_16_415 ();
 sg13g2_fill_8 FILLER_0_16_423 ();
 sg13g2_fill_4 FILLER_0_16_431 ();
 sg13g2_fill_1 FILLER_0_16_435 ();
 sg13g2_fill_2 FILLER_0_16_462 ();
 sg13g2_fill_2 FILLER_0_16_469 ();
 sg13g2_fill_8 FILLER_0_16_475 ();
 sg13g2_fill_8 FILLER_0_16_483 ();
 sg13g2_fill_8 FILLER_0_16_491 ();
 sg13g2_fill_1 FILLER_0_16_499 ();
 sg13g2_fill_2 FILLER_0_16_526 ();
 sg13g2_fill_1 FILLER_0_16_528 ();
 sg13g2_fill_8 FILLER_0_16_534 ();
 sg13g2_fill_8 FILLER_0_16_542 ();
 sg13g2_fill_4 FILLER_0_16_550 ();
 sg13g2_fill_8 FILLER_0_16_559 ();
 sg13g2_fill_8 FILLER_0_16_567 ();
 sg13g2_fill_8 FILLER_0_16_575 ();
 sg13g2_fill_8 FILLER_0_16_583 ();
 sg13g2_fill_8 FILLER_0_16_591 ();
 sg13g2_fill_1 FILLER_0_16_599 ();
 sg13g2_fill_2 FILLER_0_16_626 ();
 sg13g2_fill_2 FILLER_0_16_633 ();
 sg13g2_fill_1 FILLER_0_16_635 ();
 sg13g2_fill_8 FILLER_0_16_641 ();
 sg13g2_fill_1 FILLER_0_16_649 ();
 sg13g2_fill_8 FILLER_0_16_676 ();
 sg13g2_fill_8 FILLER_0_16_684 ();
 sg13g2_fill_1 FILLER_0_16_692 ();
 sg13g2_fill_8 FILLER_0_16_698 ();
 sg13g2_fill_8 FILLER_0_16_706 ();
 sg13g2_fill_2 FILLER_0_16_714 ();
 sg13g2_fill_8 FILLER_0_16_721 ();
 sg13g2_fill_4 FILLER_0_16_734 ();
 sg13g2_fill_4 FILLER_0_16_743 ();
 sg13g2_fill_2 FILLER_0_16_752 ();
 sg13g2_fill_1 FILLER_0_16_754 ();
 sg13g2_fill_2 FILLER_0_16_760 ();
 sg13g2_fill_2 FILLER_0_16_766 ();
 sg13g2_fill_1 FILLER_0_16_768 ();
 sg13g2_fill_2 FILLER_0_16_775 ();
 sg13g2_fill_2 FILLER_0_16_784 ();
 sg13g2_fill_2 FILLER_0_16_791 ();
 sg13g2_fill_2 FILLER_0_16_798 ();
 sg13g2_fill_2 FILLER_0_16_805 ();
 sg13g2_fill_2 FILLER_0_16_812 ();
 sg13g2_fill_2 FILLER_0_16_819 ();
 sg13g2_fill_2 FILLER_0_16_825 ();
 sg13g2_fill_2 FILLER_0_16_835 ();
 sg13g2_fill_2 FILLER_0_16_858 ();
 sg13g2_fill_1 FILLER_0_16_860 ();
 sg13g2_fill_8 FILLER_0_16_866 ();
 sg13g2_fill_4 FILLER_0_16_874 ();
 sg13g2_fill_1 FILLER_0_16_878 ();
 sg13g2_fill_2 FILLER_0_16_884 ();
 sg13g2_fill_1 FILLER_0_16_886 ();
 sg13g2_fill_2 FILLER_0_16_891 ();
 sg13g2_fill_8 FILLER_0_16_898 ();
 sg13g2_fill_4 FILLER_0_16_906 ();
 sg13g2_fill_2 FILLER_0_16_936 ();
 sg13g2_fill_2 FILLER_0_16_943 ();
 sg13g2_fill_1 FILLER_0_16_945 ();
 sg13g2_fill_8 FILLER_0_16_950 ();
 sg13g2_fill_8 FILLER_0_16_958 ();
 sg13g2_fill_8 FILLER_0_16_966 ();
 sg13g2_fill_1 FILLER_0_16_974 ();
 sg13g2_fill_2 FILLER_0_16_980 ();
 sg13g2_fill_2 FILLER_0_16_986 ();
 sg13g2_fill_4 FILLER_0_16_994 ();
 sg13g2_fill_8 FILLER_0_16_1024 ();
 sg13g2_fill_2 FILLER_0_16_1032 ();
 sg13g2_fill_8 FILLER_0_16_1040 ();
 sg13g2_fill_8 FILLER_0_16_1048 ();
 sg13g2_fill_8 FILLER_0_16_1056 ();
 sg13g2_fill_4 FILLER_0_16_1064 ();
 sg13g2_fill_2 FILLER_0_16_1068 ();
 sg13g2_fill_8 FILLER_0_16_1074 ();
 sg13g2_fill_8 FILLER_0_16_1087 ();
 sg13g2_fill_8 FILLER_0_16_1095 ();
 sg13g2_fill_8 FILLER_0_16_1103 ();
 sg13g2_fill_8 FILLER_0_16_1111 ();
 sg13g2_fill_4 FILLER_0_16_1119 ();
 sg13g2_fill_2 FILLER_0_16_1149 ();
 sg13g2_fill_8 FILLER_0_16_1172 ();
 sg13g2_fill_4 FILLER_0_16_1180 ();
 sg13g2_fill_2 FILLER_0_16_1184 ();
 sg13g2_fill_1 FILLER_0_16_1186 ();
 sg13g2_fill_2 FILLER_0_16_1213 ();
 sg13g2_fill_8 FILLER_0_16_1236 ();
 sg13g2_fill_8 FILLER_0_16_1244 ();
 sg13g2_fill_8 FILLER_0_16_1252 ();
 sg13g2_fill_8 FILLER_0_16_1260 ();
 sg13g2_fill_8 FILLER_0_16_1268 ();
 sg13g2_fill_8 FILLER_0_16_1276 ();
 sg13g2_fill_8 FILLER_0_16_1284 ();
 sg13g2_fill_4 FILLER_0_16_1292 ();
 sg13g2_fill_1 FILLER_0_16_1296 ();
 sg13g2_fill_8 FILLER_0_17_0 ();
 sg13g2_fill_8 FILLER_0_17_8 ();
 sg13g2_fill_8 FILLER_0_17_16 ();
 sg13g2_fill_8 FILLER_0_17_24 ();
 sg13g2_fill_8 FILLER_0_17_32 ();
 sg13g2_fill_8 FILLER_0_17_40 ();
 sg13g2_fill_8 FILLER_0_17_48 ();
 sg13g2_fill_8 FILLER_0_17_56 ();
 sg13g2_fill_8 FILLER_0_17_64 ();
 sg13g2_fill_8 FILLER_0_17_72 ();
 sg13g2_fill_8 FILLER_0_17_80 ();
 sg13g2_fill_8 FILLER_0_17_88 ();
 sg13g2_fill_8 FILLER_0_17_96 ();
 sg13g2_fill_8 FILLER_0_17_104 ();
 sg13g2_fill_8 FILLER_0_17_112 ();
 sg13g2_fill_8 FILLER_0_17_120 ();
 sg13g2_fill_8 FILLER_0_17_128 ();
 sg13g2_fill_8 FILLER_0_17_136 ();
 sg13g2_fill_8 FILLER_0_17_144 ();
 sg13g2_fill_8 FILLER_0_17_152 ();
 sg13g2_fill_8 FILLER_0_17_160 ();
 sg13g2_fill_8 FILLER_0_17_168 ();
 sg13g2_fill_8 FILLER_0_17_176 ();
 sg13g2_fill_8 FILLER_0_17_184 ();
 sg13g2_fill_8 FILLER_0_17_192 ();
 sg13g2_fill_8 FILLER_0_17_200 ();
 sg13g2_fill_8 FILLER_0_17_208 ();
 sg13g2_fill_8 FILLER_0_17_216 ();
 sg13g2_fill_8 FILLER_0_17_224 ();
 sg13g2_fill_8 FILLER_0_17_232 ();
 sg13g2_fill_8 FILLER_0_17_240 ();
 sg13g2_fill_8 FILLER_0_17_248 ();
 sg13g2_fill_8 FILLER_0_17_256 ();
 sg13g2_fill_8 FILLER_0_17_264 ();
 sg13g2_fill_8 FILLER_0_17_272 ();
 sg13g2_fill_8 FILLER_0_17_280 ();
 sg13g2_fill_8 FILLER_0_17_288 ();
 sg13g2_fill_2 FILLER_0_17_296 ();
 sg13g2_fill_1 FILLER_0_17_298 ();
 sg13g2_fill_2 FILLER_0_17_325 ();
 sg13g2_fill_1 FILLER_0_17_327 ();
 sg13g2_fill_4 FILLER_0_17_333 ();
 sg13g2_fill_2 FILLER_0_17_342 ();
 sg13g2_fill_8 FILLER_0_17_348 ();
 sg13g2_fill_8 FILLER_0_17_356 ();
 sg13g2_fill_8 FILLER_0_17_364 ();
 sg13g2_fill_2 FILLER_0_17_377 ();
 sg13g2_fill_2 FILLER_0_17_384 ();
 sg13g2_fill_2 FILLER_0_17_392 ();
 sg13g2_fill_1 FILLER_0_17_394 ();
 sg13g2_fill_2 FILLER_0_17_400 ();
 sg13g2_fill_1 FILLER_0_17_402 ();
 sg13g2_fill_2 FILLER_0_17_408 ();
 sg13g2_fill_4 FILLER_0_17_436 ();
 sg13g2_fill_2 FILLER_0_17_445 ();
 sg13g2_fill_2 FILLER_0_17_452 ();
 sg13g2_fill_8 FILLER_0_17_480 ();
 sg13g2_fill_8 FILLER_0_17_488 ();
 sg13g2_fill_8 FILLER_0_17_496 ();
 sg13g2_fill_8 FILLER_0_17_504 ();
 sg13g2_fill_1 FILLER_0_17_512 ();
 sg13g2_fill_2 FILLER_0_17_539 ();
 sg13g2_fill_4 FILLER_0_17_548 ();
 sg13g2_fill_8 FILLER_0_17_557 ();
 sg13g2_fill_2 FILLER_0_17_565 ();
 sg13g2_fill_1 FILLER_0_17_567 ();
 sg13g2_fill_8 FILLER_0_17_573 ();
 sg13g2_fill_4 FILLER_0_17_581 ();
 sg13g2_fill_8 FILLER_0_17_611 ();
 sg13g2_fill_4 FILLER_0_17_619 ();
 sg13g2_fill_2 FILLER_0_17_628 ();
 sg13g2_fill_8 FILLER_0_17_637 ();
 sg13g2_fill_8 FILLER_0_17_645 ();
 sg13g2_fill_2 FILLER_0_17_658 ();
 sg13g2_fill_8 FILLER_0_17_664 ();
 sg13g2_fill_4 FILLER_0_17_672 ();
 sg13g2_fill_1 FILLER_0_17_676 ();
 sg13g2_fill_4 FILLER_0_17_682 ();
 sg13g2_fill_1 FILLER_0_17_686 ();
 sg13g2_fill_8 FILLER_0_17_692 ();
 sg13g2_fill_2 FILLER_0_17_705 ();
 sg13g2_fill_2 FILLER_0_17_712 ();
 sg13g2_fill_8 FILLER_0_17_740 ();
 sg13g2_fill_4 FILLER_0_17_748 ();
 sg13g2_fill_2 FILLER_0_17_757 ();
 sg13g2_fill_1 FILLER_0_17_759 ();
 sg13g2_fill_4 FILLER_0_17_764 ();
 sg13g2_fill_1 FILLER_0_17_768 ();
 sg13g2_fill_8 FILLER_0_17_795 ();
 sg13g2_fill_4 FILLER_0_17_829 ();
 sg13g2_fill_1 FILLER_0_17_833 ();
 sg13g2_fill_8 FILLER_0_17_839 ();
 sg13g2_fill_8 FILLER_0_17_855 ();
 sg13g2_fill_2 FILLER_0_17_863 ();
 sg13g2_fill_1 FILLER_0_17_865 ();
 sg13g2_fill_2 FILLER_0_17_870 ();
 sg13g2_fill_2 FILLER_0_17_878 ();
 sg13g2_fill_2 FILLER_0_17_890 ();
 sg13g2_fill_8 FILLER_0_17_898 ();
 sg13g2_fill_4 FILLER_0_17_906 ();
 sg13g2_fill_8 FILLER_0_17_915 ();
 sg13g2_fill_8 FILLER_0_17_923 ();
 sg13g2_fill_8 FILLER_0_17_931 ();
 sg13g2_fill_1 FILLER_0_17_939 ();
 sg13g2_fill_4 FILLER_0_17_966 ();
 sg13g2_fill_2 FILLER_0_17_970 ();
 sg13g2_fill_2 FILLER_0_17_998 ();
 sg13g2_fill_4 FILLER_0_17_1010 ();
 sg13g2_fill_2 FILLER_0_17_1020 ();
 sg13g2_fill_2 FILLER_0_17_1026 ();
 sg13g2_fill_8 FILLER_0_17_1033 ();
 sg13g2_fill_8 FILLER_0_17_1041 ();
 sg13g2_fill_1 FILLER_0_17_1049 ();
 sg13g2_fill_4 FILLER_0_17_1054 ();
 sg13g2_fill_4 FILLER_0_17_1084 ();
 sg13g2_fill_1 FILLER_0_17_1088 ();
 sg13g2_fill_2 FILLER_0_17_1110 ();
 sg13g2_fill_8 FILLER_0_17_1133 ();
 sg13g2_fill_1 FILLER_0_17_1141 ();
 sg13g2_fill_4 FILLER_0_17_1146 ();
 sg13g2_fill_2 FILLER_0_17_1150 ();
 sg13g2_fill_1 FILLER_0_17_1152 ();
 sg13g2_fill_2 FILLER_0_17_1158 ();
 sg13g2_fill_2 FILLER_0_17_1186 ();
 sg13g2_fill_1 FILLER_0_17_1188 ();
 sg13g2_fill_2 FILLER_0_17_1194 ();
 sg13g2_fill_1 FILLER_0_17_1196 ();
 sg13g2_fill_2 FILLER_0_17_1201 ();
 sg13g2_fill_1 FILLER_0_17_1203 ();
 sg13g2_fill_4 FILLER_0_17_1209 ();
 sg13g2_fill_2 FILLER_0_17_1218 ();
 sg13g2_fill_8 FILLER_0_17_1246 ();
 sg13g2_fill_8 FILLER_0_17_1254 ();
 sg13g2_fill_8 FILLER_0_17_1262 ();
 sg13g2_fill_8 FILLER_0_17_1270 ();
 sg13g2_fill_8 FILLER_0_17_1278 ();
 sg13g2_fill_8 FILLER_0_17_1286 ();
 sg13g2_fill_2 FILLER_0_17_1294 ();
 sg13g2_fill_1 FILLER_0_17_1296 ();
 sg13g2_fill_8 FILLER_0_18_0 ();
 sg13g2_fill_8 FILLER_0_18_8 ();
 sg13g2_fill_8 FILLER_0_18_16 ();
 sg13g2_fill_8 FILLER_0_18_24 ();
 sg13g2_fill_8 FILLER_0_18_32 ();
 sg13g2_fill_8 FILLER_0_18_40 ();
 sg13g2_fill_8 FILLER_0_18_48 ();
 sg13g2_fill_8 FILLER_0_18_56 ();
 sg13g2_fill_8 FILLER_0_18_64 ();
 sg13g2_fill_8 FILLER_0_18_72 ();
 sg13g2_fill_8 FILLER_0_18_80 ();
 sg13g2_fill_8 FILLER_0_18_88 ();
 sg13g2_fill_8 FILLER_0_18_96 ();
 sg13g2_fill_8 FILLER_0_18_104 ();
 sg13g2_fill_8 FILLER_0_18_112 ();
 sg13g2_fill_8 FILLER_0_18_120 ();
 sg13g2_fill_8 FILLER_0_18_128 ();
 sg13g2_fill_8 FILLER_0_18_136 ();
 sg13g2_fill_8 FILLER_0_18_144 ();
 sg13g2_fill_8 FILLER_0_18_152 ();
 sg13g2_fill_8 FILLER_0_18_160 ();
 sg13g2_fill_8 FILLER_0_18_168 ();
 sg13g2_fill_8 FILLER_0_18_176 ();
 sg13g2_fill_8 FILLER_0_18_184 ();
 sg13g2_fill_8 FILLER_0_18_192 ();
 sg13g2_fill_8 FILLER_0_18_200 ();
 sg13g2_fill_8 FILLER_0_18_208 ();
 sg13g2_fill_8 FILLER_0_18_216 ();
 sg13g2_fill_8 FILLER_0_18_224 ();
 sg13g2_fill_8 FILLER_0_18_232 ();
 sg13g2_fill_8 FILLER_0_18_240 ();
 sg13g2_fill_8 FILLER_0_18_248 ();
 sg13g2_fill_8 FILLER_0_18_256 ();
 sg13g2_fill_8 FILLER_0_18_264 ();
 sg13g2_fill_8 FILLER_0_18_272 ();
 sg13g2_fill_2 FILLER_0_18_280 ();
 sg13g2_fill_1 FILLER_0_18_282 ();
 sg13g2_fill_2 FILLER_0_18_288 ();
 sg13g2_fill_8 FILLER_0_18_294 ();
 sg13g2_fill_8 FILLER_0_18_302 ();
 sg13g2_fill_8 FILLER_0_18_310 ();
 sg13g2_fill_8 FILLER_0_18_318 ();
 sg13g2_fill_1 FILLER_0_18_326 ();
 sg13g2_fill_2 FILLER_0_18_353 ();
 sg13g2_fill_1 FILLER_0_18_355 ();
 sg13g2_fill_4 FILLER_0_18_361 ();
 sg13g2_fill_1 FILLER_0_18_365 ();
 sg13g2_fill_2 FILLER_0_18_371 ();
 sg13g2_fill_1 FILLER_0_18_373 ();
 sg13g2_fill_2 FILLER_0_18_382 ();
 sg13g2_fill_8 FILLER_0_18_390 ();
 sg13g2_fill_2 FILLER_0_18_403 ();
 sg13g2_fill_4 FILLER_0_18_409 ();
 sg13g2_fill_2 FILLER_0_18_413 ();
 sg13g2_fill_4 FILLER_0_18_441 ();
 sg13g2_fill_1 FILLER_0_18_445 ();
 sg13g2_fill_2 FILLER_0_18_467 ();
 sg13g2_fill_8 FILLER_0_18_475 ();
 sg13g2_fill_8 FILLER_0_18_483 ();
 sg13g2_fill_8 FILLER_0_18_491 ();
 sg13g2_fill_8 FILLER_0_18_499 ();
 sg13g2_fill_4 FILLER_0_18_507 ();
 sg13g2_fill_2 FILLER_0_18_511 ();
 sg13g2_fill_1 FILLER_0_18_513 ();
 sg13g2_fill_2 FILLER_0_18_519 ();
 sg13g2_fill_2 FILLER_0_18_526 ();
 sg13g2_fill_2 FILLER_0_18_533 ();
 sg13g2_fill_4 FILLER_0_18_539 ();
 sg13g2_fill_8 FILLER_0_18_548 ();
 sg13g2_fill_2 FILLER_0_18_562 ();
 sg13g2_fill_2 FILLER_0_18_576 ();
 sg13g2_fill_8 FILLER_0_18_583 ();
 sg13g2_fill_2 FILLER_0_18_591 ();
 sg13g2_fill_1 FILLER_0_18_593 ();
 sg13g2_fill_4 FILLER_0_18_598 ();
 sg13g2_fill_2 FILLER_0_18_602 ();
 sg13g2_fill_4 FILLER_0_18_609 ();
 sg13g2_fill_2 FILLER_0_18_618 ();
 sg13g2_fill_2 FILLER_0_18_625 ();
 sg13g2_fill_8 FILLER_0_18_632 ();
 sg13g2_fill_8 FILLER_0_18_640 ();
 sg13g2_fill_8 FILLER_0_18_648 ();
 sg13g2_fill_2 FILLER_0_18_656 ();
 sg13g2_fill_8 FILLER_0_18_662 ();
 sg13g2_fill_1 FILLER_0_18_670 ();
 sg13g2_fill_2 FILLER_0_18_692 ();
 sg13g2_fill_1 FILLER_0_18_694 ();
 sg13g2_fill_2 FILLER_0_18_701 ();
 sg13g2_fill_2 FILLER_0_18_708 ();
 sg13g2_fill_4 FILLER_0_18_714 ();
 sg13g2_fill_1 FILLER_0_18_718 ();
 sg13g2_fill_4 FILLER_0_18_726 ();
 sg13g2_fill_1 FILLER_0_18_730 ();
 sg13g2_fill_8 FILLER_0_18_736 ();
 sg13g2_fill_8 FILLER_0_18_744 ();
 sg13g2_fill_8 FILLER_0_18_778 ();
 sg13g2_fill_8 FILLER_0_18_786 ();
 sg13g2_fill_8 FILLER_0_18_794 ();
 sg13g2_fill_4 FILLER_0_18_802 ();
 sg13g2_fill_2 FILLER_0_18_806 ();
 sg13g2_fill_1 FILLER_0_18_808 ();
 sg13g2_fill_2 FILLER_0_18_835 ();
 sg13g2_fill_4 FILLER_0_18_847 ();
 sg13g2_fill_2 FILLER_0_18_851 ();
 sg13g2_fill_2 FILLER_0_18_879 ();
 sg13g2_fill_4 FILLER_0_18_907 ();
 sg13g2_fill_2 FILLER_0_18_915 ();
 sg13g2_fill_1 FILLER_0_18_917 ();
 sg13g2_fill_2 FILLER_0_18_926 ();
 sg13g2_fill_2 FILLER_0_18_933 ();
 sg13g2_fill_1 FILLER_0_18_935 ();
 sg13g2_fill_4 FILLER_0_18_941 ();
 sg13g2_fill_2 FILLER_0_18_950 ();
 sg13g2_fill_1 FILLER_0_18_952 ();
 sg13g2_fill_4 FILLER_0_18_958 ();
 sg13g2_fill_1 FILLER_0_18_962 ();
 sg13g2_fill_8 FILLER_0_18_968 ();
 sg13g2_fill_8 FILLER_0_18_976 ();
 sg13g2_fill_2 FILLER_0_18_984 ();
 sg13g2_fill_2 FILLER_0_18_991 ();
 sg13g2_fill_4 FILLER_0_18_998 ();
 sg13g2_fill_4 FILLER_0_18_1007 ();
 sg13g2_fill_1 FILLER_0_18_1011 ();
 sg13g2_fill_4 FILLER_0_18_1017 ();
 sg13g2_fill_4 FILLER_0_18_1025 ();
 sg13g2_fill_1 FILLER_0_18_1029 ();
 sg13g2_fill_4 FILLER_0_18_1038 ();
 sg13g2_fill_1 FILLER_0_18_1042 ();
 sg13g2_fill_2 FILLER_0_18_1048 ();
 sg13g2_fill_1 FILLER_0_18_1050 ();
 sg13g2_fill_2 FILLER_0_18_1077 ();
 sg13g2_fill_1 FILLER_0_18_1079 ();
 sg13g2_fill_2 FILLER_0_18_1085 ();
 sg13g2_fill_1 FILLER_0_18_1087 ();
 sg13g2_fill_4 FILLER_0_18_1092 ();
 sg13g2_fill_8 FILLER_0_18_1122 ();
 sg13g2_fill_2 FILLER_0_18_1135 ();
 sg13g2_fill_2 FILLER_0_18_1163 ();
 sg13g2_fill_8 FILLER_0_18_1186 ();
 sg13g2_fill_1 FILLER_0_18_1194 ();
 sg13g2_fill_2 FILLER_0_18_1221 ();
 sg13g2_fill_8 FILLER_0_18_1227 ();
 sg13g2_fill_8 FILLER_0_18_1235 ();
 sg13g2_fill_8 FILLER_0_18_1243 ();
 sg13g2_fill_8 FILLER_0_18_1251 ();
 sg13g2_fill_8 FILLER_0_18_1259 ();
 sg13g2_fill_8 FILLER_0_18_1267 ();
 sg13g2_fill_8 FILLER_0_18_1275 ();
 sg13g2_fill_8 FILLER_0_18_1283 ();
 sg13g2_fill_4 FILLER_0_18_1291 ();
 sg13g2_fill_2 FILLER_0_18_1295 ();
 sg13g2_fill_8 FILLER_0_19_0 ();
 sg13g2_fill_8 FILLER_0_19_8 ();
 sg13g2_fill_8 FILLER_0_19_16 ();
 sg13g2_fill_8 FILLER_0_19_24 ();
 sg13g2_fill_8 FILLER_0_19_32 ();
 sg13g2_fill_8 FILLER_0_19_40 ();
 sg13g2_fill_8 FILLER_0_19_48 ();
 sg13g2_fill_8 FILLER_0_19_56 ();
 sg13g2_fill_8 FILLER_0_19_64 ();
 sg13g2_fill_8 FILLER_0_19_72 ();
 sg13g2_fill_8 FILLER_0_19_80 ();
 sg13g2_fill_8 FILLER_0_19_88 ();
 sg13g2_fill_8 FILLER_0_19_96 ();
 sg13g2_fill_8 FILLER_0_19_104 ();
 sg13g2_fill_8 FILLER_0_19_112 ();
 sg13g2_fill_8 FILLER_0_19_120 ();
 sg13g2_fill_8 FILLER_0_19_128 ();
 sg13g2_fill_8 FILLER_0_19_136 ();
 sg13g2_fill_8 FILLER_0_19_144 ();
 sg13g2_fill_8 FILLER_0_19_152 ();
 sg13g2_fill_8 FILLER_0_19_160 ();
 sg13g2_fill_8 FILLER_0_19_168 ();
 sg13g2_fill_8 FILLER_0_19_176 ();
 sg13g2_fill_8 FILLER_0_19_184 ();
 sg13g2_fill_8 FILLER_0_19_192 ();
 sg13g2_fill_8 FILLER_0_19_200 ();
 sg13g2_fill_8 FILLER_0_19_208 ();
 sg13g2_fill_8 FILLER_0_19_216 ();
 sg13g2_fill_8 FILLER_0_19_224 ();
 sg13g2_fill_8 FILLER_0_19_232 ();
 sg13g2_fill_8 FILLER_0_19_240 ();
 sg13g2_fill_8 FILLER_0_19_248 ();
 sg13g2_fill_8 FILLER_0_19_256 ();
 sg13g2_fill_8 FILLER_0_19_264 ();
 sg13g2_fill_8 FILLER_0_19_272 ();
 sg13g2_fill_4 FILLER_0_19_280 ();
 sg13g2_fill_2 FILLER_0_19_284 ();
 sg13g2_fill_1 FILLER_0_19_286 ();
 sg13g2_fill_8 FILLER_0_19_313 ();
 sg13g2_fill_8 FILLER_0_19_321 ();
 sg13g2_fill_8 FILLER_0_19_329 ();
 sg13g2_fill_4 FILLER_0_19_337 ();
 sg13g2_fill_8 FILLER_0_19_346 ();
 sg13g2_fill_1 FILLER_0_19_354 ();
 sg13g2_fill_8 FILLER_0_19_360 ();
 sg13g2_fill_8 FILLER_0_19_368 ();
 sg13g2_fill_4 FILLER_0_19_376 ();
 sg13g2_fill_8 FILLER_0_19_392 ();
 sg13g2_fill_4 FILLER_0_19_400 ();
 sg13g2_fill_4 FILLER_0_19_409 ();
 sg13g2_fill_1 FILLER_0_19_413 ();
 sg13g2_fill_2 FILLER_0_19_419 ();
 sg13g2_fill_2 FILLER_0_19_425 ();
 sg13g2_fill_8 FILLER_0_19_437 ();
 sg13g2_fill_8 FILLER_0_19_445 ();
 sg13g2_fill_1 FILLER_0_19_453 ();
 sg13g2_fill_8 FILLER_0_19_458 ();
 sg13g2_fill_8 FILLER_0_19_466 ();
 sg13g2_fill_8 FILLER_0_19_474 ();
 sg13g2_fill_2 FILLER_0_19_482 ();
 sg13g2_fill_1 FILLER_0_19_484 ();
 sg13g2_fill_2 FILLER_0_19_490 ();
 sg13g2_fill_8 FILLER_0_19_496 ();
 sg13g2_fill_8 FILLER_0_19_504 ();
 sg13g2_fill_8 FILLER_0_19_512 ();
 sg13g2_fill_8 FILLER_0_19_520 ();
 sg13g2_fill_8 FILLER_0_19_528 ();
 sg13g2_fill_8 FILLER_0_19_536 ();
 sg13g2_fill_8 FILLER_0_19_544 ();
 sg13g2_fill_8 FILLER_0_19_552 ();
 sg13g2_fill_8 FILLER_0_19_560 ();
 sg13g2_fill_8 FILLER_0_19_568 ();
 sg13g2_fill_8 FILLER_0_19_576 ();
 sg13g2_fill_4 FILLER_0_19_584 ();
 sg13g2_fill_2 FILLER_0_19_588 ();
 sg13g2_fill_2 FILLER_0_19_595 ();
 sg13g2_fill_4 FILLER_0_19_605 ();
 sg13g2_fill_1 FILLER_0_19_609 ();
 sg13g2_fill_8 FILLER_0_19_616 ();
 sg13g2_fill_1 FILLER_0_19_624 ();
 sg13g2_fill_2 FILLER_0_19_629 ();
 sg13g2_fill_8 FILLER_0_19_637 ();
 sg13g2_fill_8 FILLER_0_19_645 ();
 sg13g2_fill_4 FILLER_0_19_653 ();
 sg13g2_fill_8 FILLER_0_19_662 ();
 sg13g2_fill_1 FILLER_0_19_670 ();
 sg13g2_fill_2 FILLER_0_19_676 ();
 sg13g2_fill_8 FILLER_0_19_682 ();
 sg13g2_fill_8 FILLER_0_19_690 ();
 sg13g2_fill_1 FILLER_0_19_698 ();
 sg13g2_fill_8 FILLER_0_19_703 ();
 sg13g2_fill_8 FILLER_0_19_711 ();
 sg13g2_fill_8 FILLER_0_19_719 ();
 sg13g2_fill_8 FILLER_0_19_727 ();
 sg13g2_fill_8 FILLER_0_19_735 ();
 sg13g2_fill_8 FILLER_0_19_743 ();
 sg13g2_fill_8 FILLER_0_19_751 ();
 sg13g2_fill_8 FILLER_0_19_759 ();
 sg13g2_fill_8 FILLER_0_19_767 ();
 sg13g2_fill_2 FILLER_0_19_775 ();
 sg13g2_fill_1 FILLER_0_19_777 ();
 sg13g2_fill_8 FILLER_0_19_782 ();
 sg13g2_fill_8 FILLER_0_19_790 ();
 sg13g2_fill_4 FILLER_0_19_798 ();
 sg13g2_fill_1 FILLER_0_19_802 ();
 sg13g2_fill_8 FILLER_0_19_808 ();
 sg13g2_fill_4 FILLER_0_19_816 ();
 sg13g2_fill_8 FILLER_0_19_841 ();
 sg13g2_fill_8 FILLER_0_19_854 ();
 sg13g2_fill_4 FILLER_0_19_867 ();
 sg13g2_fill_2 FILLER_0_19_871 ();
 sg13g2_fill_2 FILLER_0_19_879 ();
 sg13g2_fill_2 FILLER_0_19_886 ();
 sg13g2_fill_2 FILLER_0_19_914 ();
 sg13g2_fill_2 FILLER_0_19_921 ();
 sg13g2_fill_2 FILLER_0_19_928 ();
 sg13g2_fill_2 FILLER_0_19_937 ();
 sg13g2_fill_8 FILLER_0_19_945 ();
 sg13g2_fill_4 FILLER_0_19_953 ();
 sg13g2_fill_2 FILLER_0_19_957 ();
 sg13g2_fill_8 FILLER_0_19_963 ();
 sg13g2_fill_8 FILLER_0_19_971 ();
 sg13g2_fill_8 FILLER_0_19_979 ();
 sg13g2_fill_8 FILLER_0_19_987 ();
 sg13g2_fill_2 FILLER_0_19_995 ();
 sg13g2_fill_8 FILLER_0_19_1002 ();
 sg13g2_fill_2 FILLER_0_19_1010 ();
 sg13g2_fill_1 FILLER_0_19_1012 ();
 sg13g2_fill_2 FILLER_0_19_1039 ();
 sg13g2_fill_2 FILLER_0_19_1046 ();
 sg13g2_fill_8 FILLER_0_19_1053 ();
 sg13g2_fill_8 FILLER_0_19_1061 ();
 sg13g2_fill_2 FILLER_0_19_1069 ();
 sg13g2_fill_1 FILLER_0_19_1071 ();
 sg13g2_fill_8 FILLER_0_19_1082 ();
 sg13g2_fill_1 FILLER_0_19_1090 ();
 sg13g2_fill_2 FILLER_0_19_1095 ();
 sg13g2_fill_8 FILLER_0_19_1102 ();
 sg13g2_fill_8 FILLER_0_19_1115 ();
 sg13g2_fill_8 FILLER_0_19_1123 ();
 sg13g2_fill_8 FILLER_0_19_1131 ();
 sg13g2_fill_8 FILLER_0_19_1139 ();
 sg13g2_fill_8 FILLER_0_19_1147 ();
 sg13g2_fill_8 FILLER_0_19_1155 ();
 sg13g2_fill_8 FILLER_0_19_1163 ();
 sg13g2_fill_8 FILLER_0_19_1171 ();
 sg13g2_fill_8 FILLER_0_19_1179 ();
 sg13g2_fill_8 FILLER_0_19_1187 ();
 sg13g2_fill_8 FILLER_0_19_1200 ();
 sg13g2_fill_8 FILLER_0_19_1208 ();
 sg13g2_fill_8 FILLER_0_19_1216 ();
 sg13g2_fill_8 FILLER_0_19_1224 ();
 sg13g2_fill_8 FILLER_0_19_1232 ();
 sg13g2_fill_8 FILLER_0_19_1240 ();
 sg13g2_fill_8 FILLER_0_19_1248 ();
 sg13g2_fill_8 FILLER_0_19_1256 ();
 sg13g2_fill_8 FILLER_0_19_1264 ();
 sg13g2_fill_8 FILLER_0_19_1272 ();
 sg13g2_fill_8 FILLER_0_19_1280 ();
 sg13g2_fill_8 FILLER_0_19_1288 ();
 sg13g2_fill_1 FILLER_0_19_1296 ();
 sg13g2_fill_8 FILLER_0_20_0 ();
 sg13g2_fill_8 FILLER_0_20_8 ();
 sg13g2_fill_8 FILLER_0_20_16 ();
 sg13g2_fill_8 FILLER_0_20_24 ();
 sg13g2_fill_8 FILLER_0_20_32 ();
 sg13g2_fill_8 FILLER_0_20_40 ();
 sg13g2_fill_8 FILLER_0_20_48 ();
 sg13g2_fill_8 FILLER_0_20_56 ();
 sg13g2_fill_8 FILLER_0_20_64 ();
 sg13g2_fill_8 FILLER_0_20_72 ();
 sg13g2_fill_8 FILLER_0_20_80 ();
 sg13g2_fill_8 FILLER_0_20_88 ();
 sg13g2_fill_8 FILLER_0_20_96 ();
 sg13g2_fill_8 FILLER_0_20_104 ();
 sg13g2_fill_8 FILLER_0_20_112 ();
 sg13g2_fill_8 FILLER_0_20_120 ();
 sg13g2_fill_8 FILLER_0_20_128 ();
 sg13g2_fill_8 FILLER_0_20_136 ();
 sg13g2_fill_8 FILLER_0_20_144 ();
 sg13g2_fill_8 FILLER_0_20_152 ();
 sg13g2_fill_8 FILLER_0_20_160 ();
 sg13g2_fill_8 FILLER_0_20_168 ();
 sg13g2_fill_8 FILLER_0_20_176 ();
 sg13g2_fill_8 FILLER_0_20_184 ();
 sg13g2_fill_8 FILLER_0_20_192 ();
 sg13g2_fill_8 FILLER_0_20_200 ();
 sg13g2_fill_8 FILLER_0_20_208 ();
 sg13g2_fill_8 FILLER_0_20_216 ();
 sg13g2_fill_8 FILLER_0_20_224 ();
 sg13g2_fill_8 FILLER_0_20_232 ();
 sg13g2_fill_8 FILLER_0_20_240 ();
 sg13g2_fill_8 FILLER_0_20_248 ();
 sg13g2_fill_8 FILLER_0_20_256 ();
 sg13g2_fill_8 FILLER_0_20_290 ();
 sg13g2_fill_8 FILLER_0_20_298 ();
 sg13g2_fill_8 FILLER_0_20_306 ();
 sg13g2_fill_8 FILLER_0_20_314 ();
 sg13g2_fill_8 FILLER_0_20_322 ();
 sg13g2_fill_8 FILLER_0_20_330 ();
 sg13g2_fill_8 FILLER_0_20_338 ();
 sg13g2_fill_4 FILLER_0_20_346 ();
 sg13g2_fill_1 FILLER_0_20_350 ();
 sg13g2_fill_8 FILLER_0_20_358 ();
 sg13g2_fill_4 FILLER_0_20_366 ();
 sg13g2_fill_2 FILLER_0_20_370 ();
 sg13g2_fill_1 FILLER_0_20_372 ();
 sg13g2_fill_2 FILLER_0_20_378 ();
 sg13g2_fill_8 FILLER_0_20_386 ();
 sg13g2_fill_8 FILLER_0_20_394 ();
 sg13g2_fill_8 FILLER_0_20_402 ();
 sg13g2_fill_8 FILLER_0_20_410 ();
 sg13g2_fill_8 FILLER_0_20_418 ();
 sg13g2_fill_4 FILLER_0_20_426 ();
 sg13g2_fill_2 FILLER_0_20_430 ();
 sg13g2_fill_8 FILLER_0_20_437 ();
 sg13g2_fill_8 FILLER_0_20_445 ();
 sg13g2_fill_8 FILLER_0_20_453 ();
 sg13g2_fill_4 FILLER_0_20_466 ();
 sg13g2_fill_2 FILLER_0_20_470 ();
 sg13g2_fill_1 FILLER_0_20_472 ();
 sg13g2_fill_2 FILLER_0_20_499 ();
 sg13g2_fill_4 FILLER_0_20_506 ();
 sg13g2_fill_8 FILLER_0_20_514 ();
 sg13g2_fill_8 FILLER_0_20_522 ();
 sg13g2_fill_8 FILLER_0_20_530 ();
 sg13g2_fill_4 FILLER_0_20_538 ();
 sg13g2_fill_8 FILLER_0_20_550 ();
 sg13g2_fill_8 FILLER_0_20_558 ();
 sg13g2_fill_8 FILLER_0_20_566 ();
 sg13g2_fill_8 FILLER_0_20_574 ();
 sg13g2_fill_8 FILLER_0_20_582 ();
 sg13g2_fill_8 FILLER_0_20_590 ();
 sg13g2_fill_8 FILLER_0_20_598 ();
 sg13g2_fill_8 FILLER_0_20_606 ();
 sg13g2_fill_4 FILLER_0_20_618 ();
 sg13g2_fill_2 FILLER_0_20_622 ();
 sg13g2_fill_2 FILLER_0_20_632 ();
 sg13g2_fill_1 FILLER_0_20_634 ();
 sg13g2_fill_4 FILLER_0_20_643 ();
 sg13g2_fill_2 FILLER_0_20_673 ();
 sg13g2_fill_1 FILLER_0_20_675 ();
 sg13g2_fill_4 FILLER_0_20_702 ();
 sg13g2_fill_2 FILLER_0_20_714 ();
 sg13g2_fill_4 FILLER_0_20_720 ();
 sg13g2_fill_1 FILLER_0_20_724 ();
 sg13g2_fill_8 FILLER_0_20_733 ();
 sg13g2_fill_8 FILLER_0_20_741 ();
 sg13g2_fill_2 FILLER_0_20_749 ();
 sg13g2_fill_8 FILLER_0_20_756 ();
 sg13g2_fill_1 FILLER_0_20_764 ();
 sg13g2_fill_8 FILLER_0_20_786 ();
 sg13g2_fill_8 FILLER_0_20_794 ();
 sg13g2_fill_8 FILLER_0_20_802 ();
 sg13g2_fill_8 FILLER_0_20_810 ();
 sg13g2_fill_8 FILLER_0_20_818 ();
 sg13g2_fill_8 FILLER_0_20_826 ();
 sg13g2_fill_8 FILLER_0_20_834 ();
 sg13g2_fill_4 FILLER_0_20_842 ();
 sg13g2_fill_2 FILLER_0_20_846 ();
 sg13g2_fill_1 FILLER_0_20_848 ();
 sg13g2_fill_8 FILLER_0_20_854 ();
 sg13g2_fill_8 FILLER_0_20_862 ();
 sg13g2_fill_8 FILLER_0_20_870 ();
 sg13g2_fill_8 FILLER_0_20_878 ();
 sg13g2_fill_8 FILLER_0_20_886 ();
 sg13g2_fill_8 FILLER_0_20_894 ();
 sg13g2_fill_8 FILLER_0_20_902 ();
 sg13g2_fill_8 FILLER_0_20_910 ();
 sg13g2_fill_4 FILLER_0_20_918 ();
 sg13g2_fill_1 FILLER_0_20_922 ();
 sg13g2_fill_8 FILLER_0_20_929 ();
 sg13g2_fill_8 FILLER_0_20_937 ();
 sg13g2_fill_8 FILLER_0_20_945 ();
 sg13g2_fill_8 FILLER_0_20_953 ();
 sg13g2_fill_4 FILLER_0_20_961 ();
 sg13g2_fill_2 FILLER_0_20_965 ();
 sg13g2_fill_1 FILLER_0_20_967 ();
 sg13g2_fill_8 FILLER_0_20_994 ();
 sg13g2_fill_1 FILLER_0_20_1002 ();
 sg13g2_fill_2 FILLER_0_20_1008 ();
 sg13g2_fill_4 FILLER_0_20_1015 ();
 sg13g2_fill_1 FILLER_0_20_1019 ();
 sg13g2_fill_8 FILLER_0_20_1025 ();
 sg13g2_fill_1 FILLER_0_20_1033 ();
 sg13g2_fill_8 FILLER_0_20_1039 ();
 sg13g2_fill_8 FILLER_0_20_1047 ();
 sg13g2_fill_2 FILLER_0_20_1055 ();
 sg13g2_fill_1 FILLER_0_20_1057 ();
 sg13g2_fill_8 FILLER_0_20_1064 ();
 sg13g2_fill_8 FILLER_0_20_1072 ();
 sg13g2_fill_8 FILLER_0_20_1080 ();
 sg13g2_fill_8 FILLER_0_20_1088 ();
 sg13g2_fill_8 FILLER_0_20_1096 ();
 sg13g2_fill_2 FILLER_0_20_1104 ();
 sg13g2_fill_1 FILLER_0_20_1106 ();
 sg13g2_fill_8 FILLER_0_20_1112 ();
 sg13g2_fill_8 FILLER_0_20_1120 ();
 sg13g2_fill_8 FILLER_0_20_1128 ();
 sg13g2_fill_8 FILLER_0_20_1136 ();
 sg13g2_fill_8 FILLER_0_20_1144 ();
 sg13g2_fill_8 FILLER_0_20_1152 ();
 sg13g2_fill_8 FILLER_0_20_1160 ();
 sg13g2_fill_8 FILLER_0_20_1168 ();
 sg13g2_fill_8 FILLER_0_20_1176 ();
 sg13g2_fill_8 FILLER_0_20_1184 ();
 sg13g2_fill_8 FILLER_0_20_1192 ();
 sg13g2_fill_8 FILLER_0_20_1200 ();
 sg13g2_fill_8 FILLER_0_20_1208 ();
 sg13g2_fill_8 FILLER_0_20_1216 ();
 sg13g2_fill_8 FILLER_0_20_1224 ();
 sg13g2_fill_8 FILLER_0_20_1232 ();
 sg13g2_fill_8 FILLER_0_20_1240 ();
 sg13g2_fill_8 FILLER_0_20_1248 ();
 sg13g2_fill_8 FILLER_0_20_1256 ();
 sg13g2_fill_8 FILLER_0_20_1264 ();
 sg13g2_fill_8 FILLER_0_20_1272 ();
 sg13g2_fill_8 FILLER_0_20_1280 ();
 sg13g2_fill_8 FILLER_0_20_1288 ();
 sg13g2_fill_1 FILLER_0_20_1296 ();
 sg13g2_fill_8 FILLER_0_21_0 ();
 sg13g2_fill_8 FILLER_0_21_8 ();
 sg13g2_fill_8 FILLER_0_21_16 ();
 sg13g2_fill_8 FILLER_0_21_24 ();
 sg13g2_fill_8 FILLER_0_21_32 ();
 sg13g2_fill_8 FILLER_0_21_40 ();
 sg13g2_fill_8 FILLER_0_21_48 ();
 sg13g2_fill_8 FILLER_0_21_56 ();
 sg13g2_fill_8 FILLER_0_21_64 ();
 sg13g2_fill_8 FILLER_0_21_72 ();
 sg13g2_fill_8 FILLER_0_21_80 ();
 sg13g2_fill_8 FILLER_0_21_88 ();
 sg13g2_fill_8 FILLER_0_21_96 ();
 sg13g2_fill_8 FILLER_0_21_104 ();
 sg13g2_fill_8 FILLER_0_21_112 ();
 sg13g2_fill_8 FILLER_0_21_120 ();
 sg13g2_fill_8 FILLER_0_21_128 ();
 sg13g2_fill_8 FILLER_0_21_136 ();
 sg13g2_fill_8 FILLER_0_21_144 ();
 sg13g2_fill_8 FILLER_0_21_152 ();
 sg13g2_fill_8 FILLER_0_21_160 ();
 sg13g2_fill_8 FILLER_0_21_168 ();
 sg13g2_fill_8 FILLER_0_21_176 ();
 sg13g2_fill_8 FILLER_0_21_184 ();
 sg13g2_fill_8 FILLER_0_21_192 ();
 sg13g2_fill_8 FILLER_0_21_200 ();
 sg13g2_fill_8 FILLER_0_21_208 ();
 sg13g2_fill_8 FILLER_0_21_216 ();
 sg13g2_fill_8 FILLER_0_21_224 ();
 sg13g2_fill_8 FILLER_0_21_232 ();
 sg13g2_fill_8 FILLER_0_21_240 ();
 sg13g2_fill_8 FILLER_0_21_248 ();
 sg13g2_fill_4 FILLER_0_21_256 ();
 sg13g2_fill_2 FILLER_0_21_260 ();
 sg13g2_fill_1 FILLER_0_21_262 ();
 sg13g2_fill_4 FILLER_0_21_268 ();
 sg13g2_fill_2 FILLER_0_21_272 ();
 sg13g2_fill_1 FILLER_0_21_274 ();
 sg13g2_fill_8 FILLER_0_21_279 ();
 sg13g2_fill_4 FILLER_0_21_287 ();
 sg13g2_fill_2 FILLER_0_21_291 ();
 sg13g2_fill_1 FILLER_0_21_293 ();
 sg13g2_fill_2 FILLER_0_21_299 ();
 sg13g2_fill_2 FILLER_0_21_305 ();
 sg13g2_fill_4 FILLER_0_21_328 ();
 sg13g2_fill_2 FILLER_0_21_332 ();
 sg13g2_fill_8 FILLER_0_21_341 ();
 sg13g2_fill_8 FILLER_0_21_349 ();
 sg13g2_fill_2 FILLER_0_21_357 ();
 sg13g2_fill_1 FILLER_0_21_359 ();
 sg13g2_fill_4 FILLER_0_21_368 ();
 sg13g2_fill_2 FILLER_0_21_372 ();
 sg13g2_fill_2 FILLER_0_21_379 ();
 sg13g2_fill_8 FILLER_0_21_385 ();
 sg13g2_fill_8 FILLER_0_21_393 ();
 sg13g2_fill_2 FILLER_0_21_401 ();
 sg13g2_fill_1 FILLER_0_21_403 ();
 sg13g2_fill_8 FILLER_0_21_409 ();
 sg13g2_fill_8 FILLER_0_21_417 ();
 sg13g2_fill_8 FILLER_0_21_425 ();
 sg13g2_fill_8 FILLER_0_21_433 ();
 sg13g2_fill_8 FILLER_0_21_441 ();
 sg13g2_fill_8 FILLER_0_21_449 ();
 sg13g2_fill_8 FILLER_0_21_457 ();
 sg13g2_fill_8 FILLER_0_21_465 ();
 sg13g2_fill_8 FILLER_0_21_473 ();
 sg13g2_fill_8 FILLER_0_21_481 ();
 sg13g2_fill_4 FILLER_0_21_489 ();
 sg13g2_fill_2 FILLER_0_21_519 ();
 sg13g2_fill_1 FILLER_0_21_521 ();
 sg13g2_fill_2 FILLER_0_21_526 ();
 sg13g2_fill_2 FILLER_0_21_533 ();
 sg13g2_fill_1 FILLER_0_21_535 ();
 sg13g2_fill_2 FILLER_0_21_541 ();
 sg13g2_fill_2 FILLER_0_21_548 ();
 sg13g2_fill_8 FILLER_0_21_555 ();
 sg13g2_fill_4 FILLER_0_21_563 ();
 sg13g2_fill_8 FILLER_0_21_571 ();
 sg13g2_fill_8 FILLER_0_21_579 ();
 sg13g2_fill_2 FILLER_0_21_587 ();
 sg13g2_fill_1 FILLER_0_21_589 ();
 sg13g2_fill_8 FILLER_0_21_616 ();
 sg13g2_fill_8 FILLER_0_21_624 ();
 sg13g2_fill_8 FILLER_0_21_637 ();
 sg13g2_fill_8 FILLER_0_21_645 ();
 sg13g2_fill_8 FILLER_0_21_653 ();
 sg13g2_fill_4 FILLER_0_21_661 ();
 sg13g2_fill_2 FILLER_0_21_665 ();
 sg13g2_fill_2 FILLER_0_21_671 ();
 sg13g2_fill_1 FILLER_0_21_673 ();
 sg13g2_fill_8 FILLER_0_21_682 ();
 sg13g2_fill_8 FILLER_0_21_690 ();
 sg13g2_fill_4 FILLER_0_21_698 ();
 sg13g2_fill_2 FILLER_0_21_708 ();
 sg13g2_fill_8 FILLER_0_21_714 ();
 sg13g2_fill_8 FILLER_0_21_722 ();
 sg13g2_fill_1 FILLER_0_21_730 ();
 sg13g2_fill_8 FILLER_0_21_738 ();
 sg13g2_fill_4 FILLER_0_21_746 ();
 sg13g2_fill_8 FILLER_0_21_776 ();
 sg13g2_fill_2 FILLER_0_21_784 ();
 sg13g2_fill_8 FILLER_0_21_812 ();
 sg13g2_fill_4 FILLER_0_21_820 ();
 sg13g2_fill_2 FILLER_0_21_850 ();
 sg13g2_fill_8 FILLER_0_21_857 ();
 sg13g2_fill_8 FILLER_0_21_865 ();
 sg13g2_fill_2 FILLER_0_21_873 ();
 sg13g2_fill_8 FILLER_0_21_880 ();
 sg13g2_fill_8 FILLER_0_21_893 ();
 sg13g2_fill_2 FILLER_0_21_901 ();
 sg13g2_fill_1 FILLER_0_21_903 ();
 sg13g2_fill_4 FILLER_0_21_914 ();
 sg13g2_fill_1 FILLER_0_21_918 ();
 sg13g2_fill_8 FILLER_0_21_925 ();
 sg13g2_fill_8 FILLER_0_21_933 ();
 sg13g2_fill_8 FILLER_0_21_941 ();
 sg13g2_fill_8 FILLER_0_21_949 ();
 sg13g2_fill_8 FILLER_0_21_957 ();
 sg13g2_fill_8 FILLER_0_21_965 ();
 sg13g2_fill_8 FILLER_0_21_973 ();
 sg13g2_fill_2 FILLER_0_21_986 ();
 sg13g2_fill_2 FILLER_0_21_993 ();
 sg13g2_fill_4 FILLER_0_21_1002 ();
 sg13g2_fill_2 FILLER_0_21_1010 ();
 sg13g2_fill_2 FILLER_0_21_1020 ();
 sg13g2_fill_8 FILLER_0_21_1027 ();
 sg13g2_fill_2 FILLER_0_21_1035 ();
 sg13g2_fill_4 FILLER_0_21_1063 ();
 sg13g2_fill_2 FILLER_0_21_1067 ();
 sg13g2_fill_1 FILLER_0_21_1069 ();
 sg13g2_fill_2 FILLER_0_21_1075 ();
 sg13g2_fill_1 FILLER_0_21_1077 ();
 sg13g2_fill_2 FILLER_0_21_1084 ();
 sg13g2_fill_1 FILLER_0_21_1086 ();
 sg13g2_fill_2 FILLER_0_21_1092 ();
 sg13g2_fill_2 FILLER_0_21_1099 ();
 sg13g2_fill_4 FILLER_0_21_1108 ();
 sg13g2_fill_1 FILLER_0_21_1112 ();
 sg13g2_fill_8 FILLER_0_21_1118 ();
 sg13g2_fill_8 FILLER_0_21_1126 ();
 sg13g2_fill_8 FILLER_0_21_1134 ();
 sg13g2_fill_8 FILLER_0_21_1142 ();
 sg13g2_fill_2 FILLER_0_21_1150 ();
 sg13g2_fill_8 FILLER_0_21_1157 ();
 sg13g2_fill_8 FILLER_0_21_1173 ();
 sg13g2_fill_4 FILLER_0_21_1181 ();
 sg13g2_fill_1 FILLER_0_21_1185 ();
 sg13g2_fill_4 FILLER_0_21_1193 ();
 sg13g2_fill_2 FILLER_0_21_1205 ();
 sg13g2_fill_8 FILLER_0_21_1212 ();
 sg13g2_fill_8 FILLER_0_21_1220 ();
 sg13g2_fill_8 FILLER_0_21_1228 ();
 sg13g2_fill_8 FILLER_0_21_1236 ();
 sg13g2_fill_8 FILLER_0_21_1244 ();
 sg13g2_fill_8 FILLER_0_21_1252 ();
 sg13g2_fill_8 FILLER_0_21_1260 ();
 sg13g2_fill_8 FILLER_0_21_1268 ();
 sg13g2_fill_8 FILLER_0_21_1276 ();
 sg13g2_fill_8 FILLER_0_21_1284 ();
 sg13g2_fill_4 FILLER_0_21_1292 ();
 sg13g2_fill_1 FILLER_0_21_1296 ();
 sg13g2_fill_8 FILLER_0_22_0 ();
 sg13g2_fill_8 FILLER_0_22_8 ();
 sg13g2_fill_8 FILLER_0_22_16 ();
 sg13g2_fill_8 FILLER_0_22_24 ();
 sg13g2_fill_8 FILLER_0_22_32 ();
 sg13g2_fill_8 FILLER_0_22_40 ();
 sg13g2_fill_8 FILLER_0_22_48 ();
 sg13g2_fill_8 FILLER_0_22_56 ();
 sg13g2_fill_8 FILLER_0_22_64 ();
 sg13g2_fill_8 FILLER_0_22_72 ();
 sg13g2_fill_8 FILLER_0_22_80 ();
 sg13g2_fill_8 FILLER_0_22_88 ();
 sg13g2_fill_8 FILLER_0_22_96 ();
 sg13g2_fill_8 FILLER_0_22_104 ();
 sg13g2_fill_8 FILLER_0_22_112 ();
 sg13g2_fill_8 FILLER_0_22_120 ();
 sg13g2_fill_8 FILLER_0_22_128 ();
 sg13g2_fill_8 FILLER_0_22_136 ();
 sg13g2_fill_8 FILLER_0_22_144 ();
 sg13g2_fill_8 FILLER_0_22_152 ();
 sg13g2_fill_8 FILLER_0_22_160 ();
 sg13g2_fill_8 FILLER_0_22_168 ();
 sg13g2_fill_8 FILLER_0_22_176 ();
 sg13g2_fill_8 FILLER_0_22_184 ();
 sg13g2_fill_8 FILLER_0_22_192 ();
 sg13g2_fill_8 FILLER_0_22_200 ();
 sg13g2_fill_8 FILLER_0_22_208 ();
 sg13g2_fill_8 FILLER_0_22_216 ();
 sg13g2_fill_8 FILLER_0_22_224 ();
 sg13g2_fill_8 FILLER_0_22_232 ();
 sg13g2_fill_4 FILLER_0_22_240 ();
 sg13g2_fill_1 FILLER_0_22_244 ();
 sg13g2_fill_8 FILLER_0_22_249 ();
 sg13g2_fill_8 FILLER_0_22_257 ();
 sg13g2_fill_8 FILLER_0_22_265 ();
 sg13g2_fill_8 FILLER_0_22_299 ();
 sg13g2_fill_4 FILLER_0_22_307 ();
 sg13g2_fill_8 FILLER_0_22_332 ();
 sg13g2_fill_4 FILLER_0_22_366 ();
 sg13g2_fill_2 FILLER_0_22_396 ();
 sg13g2_fill_2 FILLER_0_22_402 ();
 sg13g2_fill_8 FILLER_0_22_409 ();
 sg13g2_fill_2 FILLER_0_22_417 ();
 sg13g2_fill_1 FILLER_0_22_419 ();
 sg13g2_fill_4 FILLER_0_22_446 ();
 sg13g2_fill_8 FILLER_0_22_455 ();
 sg13g2_fill_1 FILLER_0_22_463 ();
 sg13g2_fill_4 FILLER_0_22_470 ();
 sg13g2_fill_2 FILLER_0_22_474 ();
 sg13g2_fill_2 FILLER_0_22_481 ();
 sg13g2_fill_1 FILLER_0_22_483 ();
 sg13g2_fill_4 FILLER_0_22_488 ();
 sg13g2_fill_4 FILLER_0_22_496 ();
 sg13g2_fill_2 FILLER_0_22_500 ();
 sg13g2_fill_2 FILLER_0_22_523 ();
 sg13g2_fill_1 FILLER_0_22_525 ();
 sg13g2_fill_4 FILLER_0_22_552 ();
 sg13g2_fill_4 FILLER_0_22_582 ();
 sg13g2_fill_8 FILLER_0_22_591 ();
 sg13g2_fill_8 FILLER_0_22_599 ();
 sg13g2_fill_8 FILLER_0_22_607 ();
 sg13g2_fill_8 FILLER_0_22_615 ();
 sg13g2_fill_8 FILLER_0_22_623 ();
 sg13g2_fill_8 FILLER_0_22_631 ();
 sg13g2_fill_8 FILLER_0_22_643 ();
 sg13g2_fill_8 FILLER_0_22_651 ();
 sg13g2_fill_4 FILLER_0_22_659 ();
 sg13g2_fill_8 FILLER_0_22_667 ();
 sg13g2_fill_8 FILLER_0_22_675 ();
 sg13g2_fill_4 FILLER_0_22_683 ();
 sg13g2_fill_1 FILLER_0_22_687 ();
 sg13g2_fill_2 FILLER_0_22_714 ();
 sg13g2_fill_1 FILLER_0_22_716 ();
 sg13g2_fill_8 FILLER_0_22_721 ();
 sg13g2_fill_4 FILLER_0_22_729 ();
 sg13g2_fill_2 FILLER_0_22_738 ();
 sg13g2_fill_2 FILLER_0_22_744 ();
 sg13g2_fill_2 FILLER_0_22_772 ();
 sg13g2_fill_2 FILLER_0_22_778 ();
 sg13g2_fill_1 FILLER_0_22_780 ();
 sg13g2_fill_2 FILLER_0_22_786 ();
 sg13g2_fill_8 FILLER_0_22_792 ();
 sg13g2_fill_8 FILLER_0_22_800 ();
 sg13g2_fill_2 FILLER_0_22_808 ();
 sg13g2_fill_1 FILLER_0_22_810 ();
 sg13g2_fill_2 FILLER_0_22_816 ();
 sg13g2_fill_1 FILLER_0_22_818 ();
 sg13g2_fill_8 FILLER_0_22_823 ();
 sg13g2_fill_8 FILLER_0_22_831 ();
 sg13g2_fill_4 FILLER_0_22_839 ();
 sg13g2_fill_2 FILLER_0_22_843 ();
 sg13g2_fill_1 FILLER_0_22_845 ();
 sg13g2_fill_4 FILLER_0_22_851 ();
 sg13g2_fill_8 FILLER_0_22_860 ();
 sg13g2_fill_8 FILLER_0_22_868 ();
 sg13g2_fill_8 FILLER_0_22_876 ();
 sg13g2_fill_4 FILLER_0_22_884 ();
 sg13g2_fill_2 FILLER_0_22_888 ();
 sg13g2_fill_1 FILLER_0_22_890 ();
 sg13g2_fill_8 FILLER_0_22_896 ();
 sg13g2_fill_8 FILLER_0_22_904 ();
 sg13g2_fill_1 FILLER_0_22_912 ();
 sg13g2_fill_2 FILLER_0_22_918 ();
 sg13g2_fill_2 FILLER_0_22_925 ();
 sg13g2_fill_1 FILLER_0_22_927 ();
 sg13g2_fill_8 FILLER_0_22_932 ();
 sg13g2_fill_8 FILLER_0_22_940 ();
 sg13g2_fill_8 FILLER_0_22_948 ();
 sg13g2_fill_8 FILLER_0_22_956 ();
 sg13g2_fill_4 FILLER_0_22_964 ();
 sg13g2_fill_1 FILLER_0_22_968 ();
 sg13g2_fill_4 FILLER_0_22_974 ();
 sg13g2_fill_2 FILLER_0_22_978 ();
 sg13g2_fill_2 FILLER_0_22_985 ();
 sg13g2_fill_2 FILLER_0_22_991 ();
 sg13g2_fill_8 FILLER_0_22_998 ();
 sg13g2_fill_8 FILLER_0_22_1006 ();
 sg13g2_fill_2 FILLER_0_22_1014 ();
 sg13g2_fill_2 FILLER_0_22_1021 ();
 sg13g2_fill_4 FILLER_0_22_1049 ();
 sg13g2_fill_8 FILLER_0_22_1063 ();
 sg13g2_fill_8 FILLER_0_22_1071 ();
 sg13g2_fill_4 FILLER_0_22_1079 ();
 sg13g2_fill_2 FILLER_0_22_1083 ();
 sg13g2_fill_8 FILLER_0_22_1111 ();
 sg13g2_fill_8 FILLER_0_22_1119 ();
 sg13g2_fill_4 FILLER_0_22_1127 ();
 sg13g2_fill_2 FILLER_0_22_1131 ();
 sg13g2_fill_2 FILLER_0_22_1159 ();
 sg13g2_fill_4 FILLER_0_22_1166 ();
 sg13g2_fill_2 FILLER_0_22_1196 ();
 sg13g2_fill_4 FILLER_0_22_1208 ();
 sg13g2_fill_2 FILLER_0_22_1212 ();
 sg13g2_fill_2 FILLER_0_22_1222 ();
 sg13g2_fill_8 FILLER_0_22_1250 ();
 sg13g2_fill_8 FILLER_0_22_1258 ();
 sg13g2_fill_8 FILLER_0_22_1266 ();
 sg13g2_fill_8 FILLER_0_22_1274 ();
 sg13g2_fill_8 FILLER_0_22_1282 ();
 sg13g2_fill_4 FILLER_0_22_1290 ();
 sg13g2_fill_2 FILLER_0_22_1294 ();
 sg13g2_fill_1 FILLER_0_22_1296 ();
 sg13g2_fill_8 FILLER_0_23_0 ();
 sg13g2_fill_8 FILLER_0_23_8 ();
 sg13g2_fill_8 FILLER_0_23_16 ();
 sg13g2_fill_8 FILLER_0_23_24 ();
 sg13g2_fill_8 FILLER_0_23_32 ();
 sg13g2_fill_8 FILLER_0_23_40 ();
 sg13g2_fill_8 FILLER_0_23_48 ();
 sg13g2_fill_8 FILLER_0_23_56 ();
 sg13g2_fill_8 FILLER_0_23_64 ();
 sg13g2_fill_8 FILLER_0_23_72 ();
 sg13g2_fill_8 FILLER_0_23_80 ();
 sg13g2_fill_8 FILLER_0_23_88 ();
 sg13g2_fill_8 FILLER_0_23_96 ();
 sg13g2_fill_8 FILLER_0_23_104 ();
 sg13g2_fill_8 FILLER_0_23_112 ();
 sg13g2_fill_8 FILLER_0_23_120 ();
 sg13g2_fill_8 FILLER_0_23_128 ();
 sg13g2_fill_8 FILLER_0_23_136 ();
 sg13g2_fill_8 FILLER_0_23_144 ();
 sg13g2_fill_8 FILLER_0_23_152 ();
 sg13g2_fill_8 FILLER_0_23_160 ();
 sg13g2_fill_8 FILLER_0_23_168 ();
 sg13g2_fill_8 FILLER_0_23_176 ();
 sg13g2_fill_8 FILLER_0_23_184 ();
 sg13g2_fill_8 FILLER_0_23_192 ();
 sg13g2_fill_8 FILLER_0_23_200 ();
 sg13g2_fill_8 FILLER_0_23_208 ();
 sg13g2_fill_8 FILLER_0_23_216 ();
 sg13g2_fill_8 FILLER_0_23_224 ();
 sg13g2_fill_2 FILLER_0_23_232 ();
 sg13g2_fill_1 FILLER_0_23_234 ();
 sg13g2_fill_2 FILLER_0_23_261 ();
 sg13g2_fill_4 FILLER_0_23_268 ();
 sg13g2_fill_2 FILLER_0_23_272 ();
 sg13g2_fill_2 FILLER_0_23_279 ();
 sg13g2_fill_8 FILLER_0_23_285 ();
 sg13g2_fill_2 FILLER_0_23_293 ();
 sg13g2_fill_1 FILLER_0_23_295 ();
 sg13g2_fill_8 FILLER_0_23_322 ();
 sg13g2_fill_8 FILLER_0_23_330 ();
 sg13g2_fill_4 FILLER_0_23_338 ();
 sg13g2_fill_1 FILLER_0_23_342 ();
 sg13g2_fill_2 FILLER_0_23_348 ();
 sg13g2_fill_1 FILLER_0_23_350 ();
 sg13g2_fill_4 FILLER_0_23_355 ();
 sg13g2_fill_1 FILLER_0_23_359 ();
 sg13g2_fill_2 FILLER_0_23_364 ();
 sg13g2_fill_8 FILLER_0_23_374 ();
 sg13g2_fill_4 FILLER_0_23_382 ();
 sg13g2_fill_4 FILLER_0_23_391 ();
 sg13g2_fill_4 FILLER_0_23_399 ();
 sg13g2_fill_1 FILLER_0_23_403 ();
 sg13g2_fill_4 FILLER_0_23_409 ();
 sg13g2_fill_2 FILLER_0_23_413 ();
 sg13g2_fill_1 FILLER_0_23_415 ();
 sg13g2_fill_2 FILLER_0_23_421 ();
 sg13g2_fill_2 FILLER_0_23_427 ();
 sg13g2_fill_4 FILLER_0_23_455 ();
 sg13g2_fill_2 FILLER_0_23_459 ();
 sg13g2_fill_1 FILLER_0_23_461 ();
 sg13g2_fill_4 FILLER_0_23_468 ();
 sg13g2_fill_2 FILLER_0_23_498 ();
 sg13g2_fill_2 FILLER_0_23_506 ();
 sg13g2_fill_8 FILLER_0_23_513 ();
 sg13g2_fill_8 FILLER_0_23_521 ();
 sg13g2_fill_2 FILLER_0_23_529 ();
 sg13g2_fill_2 FILLER_0_23_535 ();
 sg13g2_fill_8 FILLER_0_23_545 ();
 sg13g2_fill_8 FILLER_0_23_553 ();
 sg13g2_fill_2 FILLER_0_23_561 ();
 sg13g2_fill_2 FILLER_0_23_568 ();
 sg13g2_fill_2 FILLER_0_23_596 ();
 sg13g2_fill_4 FILLER_0_23_619 ();
 sg13g2_fill_1 FILLER_0_23_623 ();
 sg13g2_fill_8 FILLER_0_23_650 ();
 sg13g2_fill_2 FILLER_0_23_658 ();
 sg13g2_fill_4 FILLER_0_23_665 ();
 sg13g2_fill_2 FILLER_0_23_669 ();
 sg13g2_fill_1 FILLER_0_23_671 ();
 sg13g2_fill_2 FILLER_0_23_678 ();
 sg13g2_fill_2 FILLER_0_23_685 ();
 sg13g2_fill_1 FILLER_0_23_687 ();
 sg13g2_fill_8 FILLER_0_23_696 ();
 sg13g2_fill_2 FILLER_0_23_709 ();
 sg13g2_fill_2 FILLER_0_23_716 ();
 sg13g2_fill_8 FILLER_0_23_723 ();
 sg13g2_fill_8 FILLER_0_23_731 ();
 sg13g2_fill_2 FILLER_0_23_739 ();
 sg13g2_fill_1 FILLER_0_23_741 ();
 sg13g2_fill_4 FILLER_0_23_750 ();
 sg13g2_fill_4 FILLER_0_23_759 ();
 sg13g2_fill_2 FILLER_0_23_763 ();
 sg13g2_fill_8 FILLER_0_23_786 ();
 sg13g2_fill_8 FILLER_0_23_794 ();
 sg13g2_fill_2 FILLER_0_23_807 ();
 sg13g2_fill_2 FILLER_0_23_835 ();
 sg13g2_fill_2 FILLER_0_23_842 ();
 sg13g2_fill_4 FILLER_0_23_849 ();
 sg13g2_fill_2 FILLER_0_23_859 ();
 sg13g2_fill_2 FILLER_0_23_866 ();
 sg13g2_fill_2 FILLER_0_23_873 ();
 sg13g2_fill_2 FILLER_0_23_901 ();
 sg13g2_fill_2 FILLER_0_23_908 ();
 sg13g2_fill_4 FILLER_0_23_915 ();
 sg13g2_fill_1 FILLER_0_23_919 ();
 sg13g2_fill_2 FILLER_0_23_946 ();
 sg13g2_fill_4 FILLER_0_23_952 ();
 sg13g2_fill_2 FILLER_0_23_956 ();
 sg13g2_fill_2 FILLER_0_23_963 ();
 sg13g2_fill_1 FILLER_0_23_965 ();
 sg13g2_fill_8 FILLER_0_23_970 ();
 sg13g2_fill_8 FILLER_0_23_978 ();
 sg13g2_fill_8 FILLER_0_23_986 ();
 sg13g2_fill_8 FILLER_0_23_994 ();
 sg13g2_fill_8 FILLER_0_23_1002 ();
 sg13g2_fill_8 FILLER_0_23_1010 ();
 sg13g2_fill_2 FILLER_0_23_1018 ();
 sg13g2_fill_2 FILLER_0_23_1025 ();
 sg13g2_fill_4 FILLER_0_23_1031 ();
 sg13g2_fill_2 FILLER_0_23_1035 ();
 sg13g2_fill_2 FILLER_0_23_1042 ();
 sg13g2_fill_8 FILLER_0_23_1048 ();
 sg13g2_fill_8 FILLER_0_23_1056 ();
 sg13g2_fill_8 FILLER_0_23_1064 ();
 sg13g2_fill_8 FILLER_0_23_1072 ();
 sg13g2_fill_4 FILLER_0_23_1080 ();
 sg13g2_fill_1 FILLER_0_23_1084 ();
 sg13g2_fill_8 FILLER_0_23_1090 ();
 sg13g2_fill_8 FILLER_0_23_1098 ();
 sg13g2_fill_8 FILLER_0_23_1106 ();
 sg13g2_fill_8 FILLER_0_23_1114 ();
 sg13g2_fill_8 FILLER_0_23_1122 ();
 sg13g2_fill_8 FILLER_0_23_1130 ();
 sg13g2_fill_8 FILLER_0_23_1138 ();
 sg13g2_fill_2 FILLER_0_23_1154 ();
 sg13g2_fill_1 FILLER_0_23_1156 ();
 sg13g2_fill_2 FILLER_0_23_1167 ();
 sg13g2_fill_8 FILLER_0_23_1179 ();
 sg13g2_fill_8 FILLER_0_23_1187 ();
 sg13g2_fill_4 FILLER_0_23_1195 ();
 sg13g2_fill_1 FILLER_0_23_1199 ();
 sg13g2_fill_8 FILLER_0_23_1210 ();
 sg13g2_fill_1 FILLER_0_23_1218 ();
 sg13g2_fill_8 FILLER_0_23_1229 ();
 sg13g2_fill_8 FILLER_0_23_1237 ();
 sg13g2_fill_8 FILLER_0_23_1245 ();
 sg13g2_fill_8 FILLER_0_23_1253 ();
 sg13g2_fill_8 FILLER_0_23_1261 ();
 sg13g2_fill_8 FILLER_0_23_1269 ();
 sg13g2_fill_8 FILLER_0_23_1277 ();
 sg13g2_fill_8 FILLER_0_23_1285 ();
 sg13g2_fill_4 FILLER_0_23_1293 ();
 sg13g2_fill_8 FILLER_0_24_0 ();
 sg13g2_fill_8 FILLER_0_24_8 ();
 sg13g2_fill_8 FILLER_0_24_16 ();
 sg13g2_fill_8 FILLER_0_24_24 ();
 sg13g2_fill_8 FILLER_0_24_32 ();
 sg13g2_fill_8 FILLER_0_24_40 ();
 sg13g2_fill_8 FILLER_0_24_48 ();
 sg13g2_fill_8 FILLER_0_24_56 ();
 sg13g2_fill_8 FILLER_0_24_64 ();
 sg13g2_fill_8 FILLER_0_24_72 ();
 sg13g2_fill_8 FILLER_0_24_80 ();
 sg13g2_fill_8 FILLER_0_24_88 ();
 sg13g2_fill_8 FILLER_0_24_96 ();
 sg13g2_fill_8 FILLER_0_24_104 ();
 sg13g2_fill_8 FILLER_0_24_112 ();
 sg13g2_fill_8 FILLER_0_24_120 ();
 sg13g2_fill_8 FILLER_0_24_128 ();
 sg13g2_fill_8 FILLER_0_24_136 ();
 sg13g2_fill_8 FILLER_0_24_144 ();
 sg13g2_fill_8 FILLER_0_24_152 ();
 sg13g2_fill_8 FILLER_0_24_160 ();
 sg13g2_fill_8 FILLER_0_24_168 ();
 sg13g2_fill_8 FILLER_0_24_176 ();
 sg13g2_fill_8 FILLER_0_24_184 ();
 sg13g2_fill_8 FILLER_0_24_192 ();
 sg13g2_fill_8 FILLER_0_24_200 ();
 sg13g2_fill_8 FILLER_0_24_208 ();
 sg13g2_fill_8 FILLER_0_24_216 ();
 sg13g2_fill_8 FILLER_0_24_224 ();
 sg13g2_fill_8 FILLER_0_24_232 ();
 sg13g2_fill_4 FILLER_0_24_240 ();
 sg13g2_fill_8 FILLER_0_24_249 ();
 sg13g2_fill_8 FILLER_0_24_257 ();
 sg13g2_fill_8 FILLER_0_24_265 ();
 sg13g2_fill_8 FILLER_0_24_273 ();
 sg13g2_fill_8 FILLER_0_24_281 ();
 sg13g2_fill_8 FILLER_0_24_289 ();
 sg13g2_fill_8 FILLER_0_24_297 ();
 sg13g2_fill_8 FILLER_0_24_305 ();
 sg13g2_fill_8 FILLER_0_24_313 ();
 sg13g2_fill_8 FILLER_0_24_321 ();
 sg13g2_fill_8 FILLER_0_24_329 ();
 sg13g2_fill_8 FILLER_0_24_337 ();
 sg13g2_fill_8 FILLER_0_24_345 ();
 sg13g2_fill_8 FILLER_0_24_353 ();
 sg13g2_fill_4 FILLER_0_24_361 ();
 sg13g2_fill_1 FILLER_0_24_365 ();
 sg13g2_fill_8 FILLER_0_24_372 ();
 sg13g2_fill_4 FILLER_0_24_380 ();
 sg13g2_fill_2 FILLER_0_24_384 ();
 sg13g2_fill_2 FILLER_0_24_412 ();
 sg13g2_fill_4 FILLER_0_24_419 ();
 sg13g2_fill_1 FILLER_0_24_423 ();
 sg13g2_fill_4 FILLER_0_24_428 ();
 sg13g2_fill_1 FILLER_0_24_432 ();
 sg13g2_fill_8 FILLER_0_24_438 ();
 sg13g2_fill_4 FILLER_0_24_446 ();
 sg13g2_fill_2 FILLER_0_24_454 ();
 sg13g2_fill_1 FILLER_0_24_456 ();
 sg13g2_fill_8 FILLER_0_24_460 ();
 sg13g2_fill_2 FILLER_0_24_468 ();
 sg13g2_fill_8 FILLER_0_24_474 ();
 sg13g2_fill_8 FILLER_0_24_482 ();
 sg13g2_fill_8 FILLER_0_24_490 ();
 sg13g2_fill_8 FILLER_0_24_498 ();
 sg13g2_fill_8 FILLER_0_24_506 ();
 sg13g2_fill_8 FILLER_0_24_514 ();
 sg13g2_fill_1 FILLER_0_24_522 ();
 sg13g2_fill_8 FILLER_0_24_528 ();
 sg13g2_fill_8 FILLER_0_24_536 ();
 sg13g2_fill_1 FILLER_0_24_544 ();
 sg13g2_fill_2 FILLER_0_24_549 ();
 sg13g2_fill_2 FILLER_0_24_555 ();
 sg13g2_fill_2 FILLER_0_24_562 ();
 sg13g2_fill_2 FILLER_0_24_569 ();
 sg13g2_fill_4 FILLER_0_24_575 ();
 sg13g2_fill_2 FILLER_0_24_579 ();
 sg13g2_fill_8 FILLER_0_24_591 ();
 sg13g2_fill_8 FILLER_0_24_599 ();
 sg13g2_fill_2 FILLER_0_24_612 ();
 sg13g2_fill_2 FILLER_0_24_620 ();
 sg13g2_fill_2 FILLER_0_24_628 ();
 sg13g2_fill_2 FILLER_0_24_635 ();
 sg13g2_fill_2 FILLER_0_24_641 ();
 sg13g2_fill_8 FILLER_0_24_648 ();
 sg13g2_fill_2 FILLER_0_24_682 ();
 sg13g2_fill_2 FILLER_0_24_688 ();
 sg13g2_fill_2 FILLER_0_24_695 ();
 sg13g2_fill_2 FILLER_0_24_702 ();
 sg13g2_fill_1 FILLER_0_24_704 ();
 sg13g2_fill_8 FILLER_0_24_713 ();
 sg13g2_fill_8 FILLER_0_24_721 ();
 sg13g2_fill_8 FILLER_0_24_729 ();
 sg13g2_fill_8 FILLER_0_24_737 ();
 sg13g2_fill_8 FILLER_0_24_745 ();
 sg13g2_fill_8 FILLER_0_24_753 ();
 sg13g2_fill_8 FILLER_0_24_761 ();
 sg13g2_fill_4 FILLER_0_24_769 ();
 sg13g2_fill_2 FILLER_0_24_773 ();
 sg13g2_fill_8 FILLER_0_24_779 ();
 sg13g2_fill_2 FILLER_0_24_787 ();
 sg13g2_fill_1 FILLER_0_24_789 ();
 sg13g2_fill_2 FILLER_0_24_796 ();
 sg13g2_fill_8 FILLER_0_24_803 ();
 sg13g2_fill_8 FILLER_0_24_811 ();
 sg13g2_fill_8 FILLER_0_24_819 ();
 sg13g2_fill_8 FILLER_0_24_827 ();
 sg13g2_fill_2 FILLER_0_24_835 ();
 sg13g2_fill_1 FILLER_0_24_837 ();
 sg13g2_fill_4 FILLER_0_24_842 ();
 sg13g2_fill_2 FILLER_0_24_846 ();
 sg13g2_fill_1 FILLER_0_24_848 ();
 sg13g2_fill_4 FILLER_0_24_856 ();
 sg13g2_fill_2 FILLER_0_24_860 ();
 sg13g2_fill_1 FILLER_0_24_862 ();
 sg13g2_fill_2 FILLER_0_24_868 ();
 sg13g2_fill_2 FILLER_0_24_874 ();
 sg13g2_fill_1 FILLER_0_24_876 ();
 sg13g2_fill_8 FILLER_0_24_881 ();
 sg13g2_fill_8 FILLER_0_24_889 ();
 sg13g2_fill_8 FILLER_0_24_897 ();
 sg13g2_fill_8 FILLER_0_24_905 ();
 sg13g2_fill_8 FILLER_0_24_913 ();
 sg13g2_fill_8 FILLER_0_24_921 ();
 sg13g2_fill_8 FILLER_0_24_929 ();
 sg13g2_fill_8 FILLER_0_24_937 ();
 sg13g2_fill_8 FILLER_0_24_945 ();
 sg13g2_fill_2 FILLER_0_24_953 ();
 sg13g2_fill_1 FILLER_0_24_955 ();
 sg13g2_fill_8 FILLER_0_24_982 ();
 sg13g2_fill_8 FILLER_0_24_990 ();
 sg13g2_fill_8 FILLER_0_24_998 ();
 sg13g2_fill_1 FILLER_0_24_1006 ();
 sg13g2_fill_2 FILLER_0_24_1011 ();
 sg13g2_fill_1 FILLER_0_24_1013 ();
 sg13g2_fill_4 FILLER_0_24_1021 ();
 sg13g2_fill_1 FILLER_0_24_1025 ();
 sg13g2_fill_4 FILLER_0_24_1031 ();
 sg13g2_fill_1 FILLER_0_24_1035 ();
 sg13g2_fill_8 FILLER_0_24_1057 ();
 sg13g2_fill_8 FILLER_0_24_1065 ();
 sg13g2_fill_8 FILLER_0_24_1073 ();
 sg13g2_fill_8 FILLER_0_24_1081 ();
 sg13g2_fill_8 FILLER_0_24_1089 ();
 sg13g2_fill_8 FILLER_0_24_1097 ();
 sg13g2_fill_8 FILLER_0_24_1105 ();
 sg13g2_fill_8 FILLER_0_24_1113 ();
 sg13g2_fill_2 FILLER_0_24_1121 ();
 sg13g2_fill_2 FILLER_0_24_1149 ();
 sg13g2_fill_8 FILLER_0_24_1161 ();
 sg13g2_fill_4 FILLER_0_24_1169 ();
 sg13g2_fill_8 FILLER_0_24_1181 ();
 sg13g2_fill_4 FILLER_0_24_1189 ();
 sg13g2_fill_1 FILLER_0_24_1193 ();
 sg13g2_fill_8 FILLER_0_24_1199 ();
 sg13g2_fill_2 FILLER_0_24_1212 ();
 sg13g2_fill_2 FILLER_0_24_1224 ();
 sg13g2_fill_8 FILLER_0_24_1231 ();
 sg13g2_fill_8 FILLER_0_24_1239 ();
 sg13g2_fill_8 FILLER_0_24_1247 ();
 sg13g2_fill_8 FILLER_0_24_1255 ();
 sg13g2_fill_8 FILLER_0_24_1263 ();
 sg13g2_fill_8 FILLER_0_24_1271 ();
 sg13g2_fill_8 FILLER_0_24_1279 ();
 sg13g2_fill_8 FILLER_0_24_1287 ();
 sg13g2_fill_2 FILLER_0_24_1295 ();
 sg13g2_fill_8 FILLER_0_25_0 ();
 sg13g2_fill_8 FILLER_0_25_8 ();
 sg13g2_fill_8 FILLER_0_25_16 ();
 sg13g2_fill_8 FILLER_0_25_24 ();
 sg13g2_fill_8 FILLER_0_25_32 ();
 sg13g2_fill_8 FILLER_0_25_40 ();
 sg13g2_fill_8 FILLER_0_25_48 ();
 sg13g2_fill_8 FILLER_0_25_56 ();
 sg13g2_fill_8 FILLER_0_25_64 ();
 sg13g2_fill_8 FILLER_0_25_72 ();
 sg13g2_fill_8 FILLER_0_25_80 ();
 sg13g2_fill_8 FILLER_0_25_88 ();
 sg13g2_fill_8 FILLER_0_25_96 ();
 sg13g2_fill_8 FILLER_0_25_104 ();
 sg13g2_fill_8 FILLER_0_25_112 ();
 sg13g2_fill_8 FILLER_0_25_120 ();
 sg13g2_fill_8 FILLER_0_25_128 ();
 sg13g2_fill_8 FILLER_0_25_136 ();
 sg13g2_fill_8 FILLER_0_25_144 ();
 sg13g2_fill_8 FILLER_0_25_152 ();
 sg13g2_fill_8 FILLER_0_25_160 ();
 sg13g2_fill_8 FILLER_0_25_168 ();
 sg13g2_fill_8 FILLER_0_25_176 ();
 sg13g2_fill_8 FILLER_0_25_184 ();
 sg13g2_fill_8 FILLER_0_25_192 ();
 sg13g2_fill_8 FILLER_0_25_200 ();
 sg13g2_fill_8 FILLER_0_25_208 ();
 sg13g2_fill_8 FILLER_0_25_216 ();
 sg13g2_fill_4 FILLER_0_25_224 ();
 sg13g2_fill_2 FILLER_0_25_228 ();
 sg13g2_fill_1 FILLER_0_25_230 ();
 sg13g2_fill_2 FILLER_0_25_257 ();
 sg13g2_fill_8 FILLER_0_25_264 ();
 sg13g2_fill_8 FILLER_0_25_272 ();
 sg13g2_fill_8 FILLER_0_25_280 ();
 sg13g2_fill_8 FILLER_0_25_288 ();
 sg13g2_fill_8 FILLER_0_25_296 ();
 sg13g2_fill_8 FILLER_0_25_304 ();
 sg13g2_fill_2 FILLER_0_25_317 ();
 sg13g2_fill_8 FILLER_0_25_323 ();
 sg13g2_fill_2 FILLER_0_25_331 ();
 sg13g2_fill_1 FILLER_0_25_333 ();
 sg13g2_fill_8 FILLER_0_25_339 ();
 sg13g2_fill_8 FILLER_0_25_347 ();
 sg13g2_fill_2 FILLER_0_25_363 ();
 sg13g2_fill_2 FILLER_0_25_370 ();
 sg13g2_fill_1 FILLER_0_25_372 ();
 sg13g2_fill_2 FILLER_0_25_378 ();
 sg13g2_fill_4 FILLER_0_25_385 ();
 sg13g2_fill_2 FILLER_0_25_394 ();
 sg13g2_fill_1 FILLER_0_25_396 ();
 sg13g2_fill_4 FILLER_0_25_407 ();
 sg13g2_fill_1 FILLER_0_25_411 ();
 sg13g2_fill_8 FILLER_0_25_416 ();
 sg13g2_fill_8 FILLER_0_25_424 ();
 sg13g2_fill_2 FILLER_0_25_432 ();
 sg13g2_fill_4 FILLER_0_25_439 ();
 sg13g2_fill_2 FILLER_0_25_443 ();
 sg13g2_fill_8 FILLER_0_25_449 ();
 sg13g2_fill_8 FILLER_0_25_457 ();
 sg13g2_fill_8 FILLER_0_25_465 ();
 sg13g2_fill_8 FILLER_0_25_473 ();
 sg13g2_fill_8 FILLER_0_25_481 ();
 sg13g2_fill_8 FILLER_0_25_489 ();
 sg13g2_fill_8 FILLER_0_25_497 ();
 sg13g2_fill_8 FILLER_0_25_505 ();
 sg13g2_fill_2 FILLER_0_25_539 ();
 sg13g2_fill_1 FILLER_0_25_541 ();
 sg13g2_fill_8 FILLER_0_25_563 ();
 sg13g2_fill_8 FILLER_0_25_571 ();
 sg13g2_fill_8 FILLER_0_25_579 ();
 sg13g2_fill_8 FILLER_0_25_587 ();
 sg13g2_fill_8 FILLER_0_25_595 ();
 sg13g2_fill_8 FILLER_0_25_603 ();
 sg13g2_fill_8 FILLER_0_25_611 ();
 sg13g2_fill_8 FILLER_0_25_624 ();
 sg13g2_fill_8 FILLER_0_25_632 ();
 sg13g2_fill_8 FILLER_0_25_640 ();
 sg13g2_fill_8 FILLER_0_25_648 ();
 sg13g2_fill_8 FILLER_0_25_656 ();
 sg13g2_fill_8 FILLER_0_25_664 ();
 sg13g2_fill_8 FILLER_0_25_672 ();
 sg13g2_fill_1 FILLER_0_25_680 ();
 sg13g2_fill_8 FILLER_0_25_686 ();
 sg13g2_fill_8 FILLER_0_25_694 ();
 sg13g2_fill_8 FILLER_0_25_702 ();
 sg13g2_fill_2 FILLER_0_25_710 ();
 sg13g2_fill_1 FILLER_0_25_712 ();
 sg13g2_fill_8 FILLER_0_25_718 ();
 sg13g2_fill_8 FILLER_0_25_726 ();
 sg13g2_fill_8 FILLER_0_25_734 ();
 sg13g2_fill_8 FILLER_0_25_742 ();
 sg13g2_fill_8 FILLER_0_25_750 ();
 sg13g2_fill_8 FILLER_0_25_758 ();
 sg13g2_fill_8 FILLER_0_25_766 ();
 sg13g2_fill_4 FILLER_0_25_774 ();
 sg13g2_fill_8 FILLER_0_25_782 ();
 sg13g2_fill_8 FILLER_0_25_790 ();
 sg13g2_fill_8 FILLER_0_25_798 ();
 sg13g2_fill_8 FILLER_0_25_806 ();
 sg13g2_fill_8 FILLER_0_25_814 ();
 sg13g2_fill_8 FILLER_0_25_822 ();
 sg13g2_fill_8 FILLER_0_25_830 ();
 sg13g2_fill_8 FILLER_0_25_838 ();
 sg13g2_fill_8 FILLER_0_25_846 ();
 sg13g2_fill_8 FILLER_0_25_854 ();
 sg13g2_fill_8 FILLER_0_25_862 ();
 sg13g2_fill_8 FILLER_0_25_870 ();
 sg13g2_fill_8 FILLER_0_25_878 ();
 sg13g2_fill_8 FILLER_0_25_886 ();
 sg13g2_fill_8 FILLER_0_25_894 ();
 sg13g2_fill_8 FILLER_0_25_902 ();
 sg13g2_fill_8 FILLER_0_25_910 ();
 sg13g2_fill_4 FILLER_0_25_918 ();
 sg13g2_fill_8 FILLER_0_25_927 ();
 sg13g2_fill_4 FILLER_0_25_935 ();
 sg13g2_fill_2 FILLER_0_25_939 ();
 sg13g2_fill_8 FILLER_0_25_947 ();
 sg13g2_fill_4 FILLER_0_25_955 ();
 sg13g2_fill_1 FILLER_0_25_959 ();
 sg13g2_fill_8 FILLER_0_25_970 ();
 sg13g2_fill_8 FILLER_0_25_978 ();
 sg13g2_fill_8 FILLER_0_25_986 ();
 sg13g2_fill_2 FILLER_0_25_998 ();
 sg13g2_fill_2 FILLER_0_25_1005 ();
 sg13g2_fill_8 FILLER_0_25_1033 ();
 sg13g2_fill_4 FILLER_0_25_1041 ();
 sg13g2_fill_2 FILLER_0_25_1045 ();
 sg13g2_fill_1 FILLER_0_25_1047 ();
 sg13g2_fill_2 FILLER_0_25_1053 ();
 sg13g2_fill_8 FILLER_0_25_1062 ();
 sg13g2_fill_8 FILLER_0_25_1070 ();
 sg13g2_fill_4 FILLER_0_25_1078 ();
 sg13g2_fill_8 FILLER_0_25_1087 ();
 sg13g2_fill_2 FILLER_0_25_1095 ();
 sg13g2_fill_8 FILLER_0_25_1101 ();
 sg13g2_fill_8 FILLER_0_25_1109 ();
 sg13g2_fill_8 FILLER_0_25_1117 ();
 sg13g2_fill_8 FILLER_0_25_1125 ();
 sg13g2_fill_8 FILLER_0_25_1133 ();
 sg13g2_fill_4 FILLER_0_25_1141 ();
 sg13g2_fill_2 FILLER_0_25_1145 ();
 sg13g2_fill_8 FILLER_0_25_1157 ();
 sg13g2_fill_2 FILLER_0_25_1165 ();
 sg13g2_fill_1 FILLER_0_25_1167 ();
 sg13g2_fill_8 FILLER_0_25_1176 ();
 sg13g2_fill_4 FILLER_0_25_1184 ();
 sg13g2_fill_8 FILLER_0_25_1192 ();
 sg13g2_fill_4 FILLER_0_25_1200 ();
 sg13g2_fill_1 FILLER_0_25_1204 ();
 sg13g2_fill_8 FILLER_0_25_1209 ();
 sg13g2_fill_8 FILLER_0_25_1217 ();
 sg13g2_fill_8 FILLER_0_25_1225 ();
 sg13g2_fill_8 FILLER_0_25_1233 ();
 sg13g2_fill_8 FILLER_0_25_1241 ();
 sg13g2_fill_8 FILLER_0_25_1249 ();
 sg13g2_fill_8 FILLER_0_25_1257 ();
 sg13g2_fill_8 FILLER_0_25_1265 ();
 sg13g2_fill_8 FILLER_0_25_1273 ();
 sg13g2_fill_8 FILLER_0_25_1281 ();
 sg13g2_fill_8 FILLER_0_25_1289 ();
 sg13g2_fill_8 FILLER_0_26_0 ();
 sg13g2_fill_8 FILLER_0_26_8 ();
 sg13g2_fill_8 FILLER_0_26_16 ();
 sg13g2_fill_8 FILLER_0_26_24 ();
 sg13g2_fill_8 FILLER_0_26_32 ();
 sg13g2_fill_8 FILLER_0_26_40 ();
 sg13g2_fill_8 FILLER_0_26_48 ();
 sg13g2_fill_8 FILLER_0_26_56 ();
 sg13g2_fill_8 FILLER_0_26_64 ();
 sg13g2_fill_8 FILLER_0_26_72 ();
 sg13g2_fill_8 FILLER_0_26_80 ();
 sg13g2_fill_8 FILLER_0_26_88 ();
 sg13g2_fill_8 FILLER_0_26_96 ();
 sg13g2_fill_8 FILLER_0_26_104 ();
 sg13g2_fill_8 FILLER_0_26_112 ();
 sg13g2_fill_8 FILLER_0_26_120 ();
 sg13g2_fill_8 FILLER_0_26_128 ();
 sg13g2_fill_8 FILLER_0_26_136 ();
 sg13g2_fill_8 FILLER_0_26_144 ();
 sg13g2_fill_8 FILLER_0_26_152 ();
 sg13g2_fill_8 FILLER_0_26_160 ();
 sg13g2_fill_8 FILLER_0_26_168 ();
 sg13g2_fill_8 FILLER_0_26_176 ();
 sg13g2_fill_8 FILLER_0_26_184 ();
 sg13g2_fill_8 FILLER_0_26_192 ();
 sg13g2_fill_8 FILLER_0_26_200 ();
 sg13g2_fill_8 FILLER_0_26_208 ();
 sg13g2_fill_8 FILLER_0_26_216 ();
 sg13g2_fill_4 FILLER_0_26_224 ();
 sg13g2_fill_1 FILLER_0_26_228 ();
 sg13g2_fill_2 FILLER_0_26_234 ();
 sg13g2_fill_8 FILLER_0_26_240 ();
 sg13g2_fill_2 FILLER_0_26_248 ();
 sg13g2_fill_4 FILLER_0_26_276 ();
 sg13g2_fill_2 FILLER_0_26_280 ();
 sg13g2_fill_1 FILLER_0_26_282 ();
 sg13g2_fill_2 FILLER_0_26_309 ();
 sg13g2_fill_1 FILLER_0_26_311 ();
 sg13g2_fill_4 FILLER_0_26_338 ();
 sg13g2_fill_2 FILLER_0_26_342 ();
 sg13g2_fill_2 FILLER_0_26_349 ();
 sg13g2_fill_2 FILLER_0_26_355 ();
 sg13g2_fill_8 FILLER_0_26_362 ();
 sg13g2_fill_1 FILLER_0_26_370 ();
 sg13g2_fill_2 FILLER_0_26_376 ();
 sg13g2_fill_8 FILLER_0_26_382 ();
 sg13g2_fill_8 FILLER_0_26_390 ();
 sg13g2_fill_2 FILLER_0_26_398 ();
 sg13g2_fill_1 FILLER_0_26_400 ();
 sg13g2_fill_8 FILLER_0_26_406 ();
 sg13g2_fill_8 FILLER_0_26_414 ();
 sg13g2_fill_8 FILLER_0_26_422 ();
 sg13g2_fill_8 FILLER_0_26_430 ();
 sg13g2_fill_1 FILLER_0_26_438 ();
 sg13g2_fill_2 FILLER_0_26_460 ();
 sg13g2_fill_1 FILLER_0_26_462 ();
 sg13g2_fill_2 FILLER_0_26_467 ();
 sg13g2_fill_8 FILLER_0_26_474 ();
 sg13g2_fill_8 FILLER_0_26_482 ();
 sg13g2_fill_4 FILLER_0_26_490 ();
 sg13g2_fill_2 FILLER_0_26_499 ();
 sg13g2_fill_4 FILLER_0_26_505 ();
 sg13g2_fill_4 FILLER_0_26_514 ();
 sg13g2_fill_1 FILLER_0_26_518 ();
 sg13g2_fill_4 FILLER_0_26_523 ();
 sg13g2_fill_1 FILLER_0_26_527 ();
 sg13g2_fill_8 FILLER_0_26_554 ();
 sg13g2_fill_4 FILLER_0_26_562 ();
 sg13g2_fill_2 FILLER_0_26_566 ();
 sg13g2_fill_2 FILLER_0_26_594 ();
 sg13g2_fill_8 FILLER_0_26_622 ();
 sg13g2_fill_1 FILLER_0_26_630 ();
 sg13g2_fill_2 FILLER_0_26_637 ();
 sg13g2_fill_2 FILLER_0_26_643 ();
 sg13g2_fill_8 FILLER_0_26_651 ();
 sg13g2_fill_8 FILLER_0_26_659 ();
 sg13g2_fill_8 FILLER_0_26_667 ();
 sg13g2_fill_8 FILLER_0_26_675 ();
 sg13g2_fill_8 FILLER_0_26_683 ();
 sg13g2_fill_8 FILLER_0_26_691 ();
 sg13g2_fill_8 FILLER_0_26_699 ();
 sg13g2_fill_8 FILLER_0_26_707 ();
 sg13g2_fill_8 FILLER_0_26_715 ();
 sg13g2_fill_8 FILLER_0_26_723 ();
 sg13g2_fill_4 FILLER_0_26_731 ();
 sg13g2_fill_2 FILLER_0_26_735 ();
 sg13g2_fill_1 FILLER_0_26_737 ();
 sg13g2_fill_8 FILLER_0_26_743 ();
 sg13g2_fill_4 FILLER_0_26_751 ();
 sg13g2_fill_1 FILLER_0_26_755 ();
 sg13g2_fill_8 FILLER_0_26_760 ();
 sg13g2_fill_4 FILLER_0_26_768 ();
 sg13g2_fill_2 FILLER_0_26_772 ();
 sg13g2_fill_4 FILLER_0_26_779 ();
 sg13g2_fill_2 FILLER_0_26_783 ();
 sg13g2_fill_1 FILLER_0_26_785 ();
 sg13g2_fill_8 FILLER_0_26_812 ();
 sg13g2_fill_2 FILLER_0_26_820 ();
 sg13g2_fill_1 FILLER_0_26_822 ();
 sg13g2_fill_4 FILLER_0_26_828 ();
 sg13g2_fill_2 FILLER_0_26_832 ();
 sg13g2_fill_1 FILLER_0_26_834 ();
 sg13g2_fill_8 FILLER_0_26_839 ();
 sg13g2_fill_8 FILLER_0_26_847 ();
 sg13g2_fill_4 FILLER_0_26_855 ();
 sg13g2_fill_8 FILLER_0_26_867 ();
 sg13g2_fill_8 FILLER_0_26_875 ();
 sg13g2_fill_1 FILLER_0_26_883 ();
 sg13g2_fill_2 FILLER_0_26_888 ();
 sg13g2_fill_2 FILLER_0_26_895 ();
 sg13g2_fill_2 FILLER_0_26_923 ();
 sg13g2_fill_8 FILLER_0_26_929 ();
 sg13g2_fill_2 FILLER_0_26_937 ();
 sg13g2_fill_1 FILLER_0_26_939 ();
 sg13g2_fill_4 FILLER_0_26_945 ();
 sg13g2_fill_2 FILLER_0_26_949 ();
 sg13g2_fill_2 FILLER_0_26_957 ();
 sg13g2_fill_1 FILLER_0_26_959 ();
 sg13g2_fill_2 FILLER_0_26_966 ();
 sg13g2_fill_4 FILLER_0_26_973 ();
 sg13g2_fill_2 FILLER_0_26_977 ();
 sg13g2_fill_8 FILLER_0_26_991 ();
 sg13g2_fill_4 FILLER_0_26_999 ();
 sg13g2_fill_2 FILLER_0_26_1003 ();
 sg13g2_fill_2 FILLER_0_26_1009 ();
 sg13g2_fill_2 FILLER_0_26_1037 ();
 sg13g2_fill_2 FILLER_0_26_1044 ();
 sg13g2_fill_4 FILLER_0_26_1049 ();
 sg13g2_fill_1 FILLER_0_26_1053 ();
 sg13g2_fill_8 FILLER_0_26_1059 ();
 sg13g2_fill_8 FILLER_0_26_1067 ();
 sg13g2_fill_2 FILLER_0_26_1083 ();
 sg13g2_fill_8 FILLER_0_26_1111 ();
 sg13g2_fill_8 FILLER_0_26_1119 ();
 sg13g2_fill_4 FILLER_0_26_1127 ();
 sg13g2_fill_2 FILLER_0_26_1131 ();
 sg13g2_fill_4 FILLER_0_26_1138 ();
 sg13g2_fill_2 FILLER_0_26_1142 ();
 sg13g2_fill_8 FILLER_0_26_1148 ();
 sg13g2_fill_2 FILLER_0_26_1164 ();
 sg13g2_fill_1 FILLER_0_26_1166 ();
 sg13g2_fill_4 FILLER_0_26_1175 ();
 sg13g2_fill_2 FILLER_0_26_1179 ();
 sg13g2_fill_1 FILLER_0_26_1181 ();
 sg13g2_fill_2 FILLER_0_26_1187 ();
 sg13g2_fill_2 FILLER_0_26_1194 ();
 sg13g2_fill_1 FILLER_0_26_1196 ();
 sg13g2_fill_2 FILLER_0_26_1202 ();
 sg13g2_fill_1 FILLER_0_26_1204 ();
 sg13g2_fill_2 FILLER_0_26_1209 ();
 sg13g2_fill_1 FILLER_0_26_1211 ();
 sg13g2_fill_2 FILLER_0_26_1220 ();
 sg13g2_fill_1 FILLER_0_26_1222 ();
 sg13g2_fill_8 FILLER_0_26_1226 ();
 sg13g2_fill_8 FILLER_0_26_1234 ();
 sg13g2_fill_2 FILLER_0_26_1242 ();
 sg13g2_fill_2 FILLER_0_26_1254 ();
 sg13g2_fill_8 FILLER_0_26_1282 ();
 sg13g2_fill_4 FILLER_0_26_1290 ();
 sg13g2_fill_2 FILLER_0_26_1294 ();
 sg13g2_fill_1 FILLER_0_26_1296 ();
 sg13g2_fill_8 FILLER_0_27_0 ();
 sg13g2_fill_8 FILLER_0_27_8 ();
 sg13g2_fill_8 FILLER_0_27_16 ();
 sg13g2_fill_8 FILLER_0_27_24 ();
 sg13g2_fill_8 FILLER_0_27_32 ();
 sg13g2_fill_8 FILLER_0_27_40 ();
 sg13g2_fill_8 FILLER_0_27_48 ();
 sg13g2_fill_8 FILLER_0_27_56 ();
 sg13g2_fill_8 FILLER_0_27_64 ();
 sg13g2_fill_8 FILLER_0_27_72 ();
 sg13g2_fill_8 FILLER_0_27_80 ();
 sg13g2_fill_8 FILLER_0_27_88 ();
 sg13g2_fill_8 FILLER_0_27_96 ();
 sg13g2_fill_8 FILLER_0_27_104 ();
 sg13g2_fill_8 FILLER_0_27_112 ();
 sg13g2_fill_8 FILLER_0_27_120 ();
 sg13g2_fill_8 FILLER_0_27_128 ();
 sg13g2_fill_8 FILLER_0_27_136 ();
 sg13g2_fill_8 FILLER_0_27_144 ();
 sg13g2_fill_8 FILLER_0_27_152 ();
 sg13g2_fill_8 FILLER_0_27_160 ();
 sg13g2_fill_8 FILLER_0_27_168 ();
 sg13g2_fill_8 FILLER_0_27_176 ();
 sg13g2_fill_8 FILLER_0_27_184 ();
 sg13g2_fill_8 FILLER_0_27_192 ();
 sg13g2_fill_8 FILLER_0_27_200 ();
 sg13g2_fill_8 FILLER_0_27_208 ();
 sg13g2_fill_4 FILLER_0_27_216 ();
 sg13g2_fill_2 FILLER_0_27_220 ();
 sg13g2_fill_2 FILLER_0_27_248 ();
 sg13g2_fill_4 FILLER_0_27_271 ();
 sg13g2_fill_2 FILLER_0_27_275 ();
 sg13g2_fill_1 FILLER_0_27_277 ();
 sg13g2_fill_2 FILLER_0_27_282 ();
 sg13g2_fill_1 FILLER_0_27_284 ();
 sg13g2_fill_2 FILLER_0_27_290 ();
 sg13g2_fill_4 FILLER_0_27_296 ();
 sg13g2_fill_2 FILLER_0_27_300 ();
 sg13g2_fill_8 FILLER_0_27_328 ();
 sg13g2_fill_1 FILLER_0_27_336 ();
 sg13g2_fill_4 FILLER_0_27_358 ();
 sg13g2_fill_2 FILLER_0_27_362 ();
 sg13g2_fill_1 FILLER_0_27_364 ();
 sg13g2_fill_4 FILLER_0_27_369 ();
 sg13g2_fill_8 FILLER_0_27_399 ();
 sg13g2_fill_4 FILLER_0_27_407 ();
 sg13g2_fill_1 FILLER_0_27_411 ();
 sg13g2_fill_8 FILLER_0_27_417 ();
 sg13g2_fill_2 FILLER_0_27_451 ();
 sg13g2_fill_8 FILLER_0_27_459 ();
 sg13g2_fill_8 FILLER_0_27_467 ();
 sg13g2_fill_2 FILLER_0_27_475 ();
 sg13g2_fill_1 FILLER_0_27_477 ();
 sg13g2_fill_8 FILLER_0_27_504 ();
 sg13g2_fill_8 FILLER_0_27_512 ();
 sg13g2_fill_2 FILLER_0_27_525 ();
 sg13g2_fill_4 FILLER_0_27_531 ();
 sg13g2_fill_2 FILLER_0_27_535 ();
 sg13g2_fill_8 FILLER_0_27_547 ();
 sg13g2_fill_1 FILLER_0_27_555 ();
 sg13g2_fill_2 FILLER_0_27_560 ();
 sg13g2_fill_4 FILLER_0_27_567 ();
 sg13g2_fill_8 FILLER_0_27_575 ();
 sg13g2_fill_8 FILLER_0_27_583 ();
 sg13g2_fill_2 FILLER_0_27_591 ();
 sg13g2_fill_1 FILLER_0_27_593 ();
 sg13g2_fill_2 FILLER_0_27_599 ();
 sg13g2_fill_4 FILLER_0_27_606 ();
 sg13g2_fill_2 FILLER_0_27_614 ();
 sg13g2_fill_2 FILLER_0_27_619 ();
 sg13g2_fill_2 FILLER_0_27_627 ();
 sg13g2_fill_8 FILLER_0_27_655 ();
 sg13g2_fill_2 FILLER_0_27_663 ();
 sg13g2_fill_2 FILLER_0_27_669 ();
 sg13g2_fill_2 FILLER_0_27_697 ();
 sg13g2_fill_1 FILLER_0_27_699 ();
 sg13g2_fill_4 FILLER_0_27_721 ();
 sg13g2_fill_4 FILLER_0_27_730 ();
 sg13g2_fill_4 FILLER_0_27_760 ();
 sg13g2_fill_2 FILLER_0_27_769 ();
 sg13g2_fill_1 FILLER_0_27_771 ();
 sg13g2_fill_2 FILLER_0_27_798 ();
 sg13g2_fill_2 FILLER_0_27_805 ();
 sg13g2_fill_8 FILLER_0_27_811 ();
 sg13g2_fill_2 FILLER_0_27_819 ();
 sg13g2_fill_2 FILLER_0_27_847 ();
 sg13g2_fill_8 FILLER_0_27_853 ();
 sg13g2_fill_8 FILLER_0_27_866 ();
 sg13g2_fill_8 FILLER_0_27_874 ();
 sg13g2_fill_8 FILLER_0_27_882 ();
 sg13g2_fill_4 FILLER_0_27_890 ();
 sg13g2_fill_2 FILLER_0_27_894 ();
 sg13g2_fill_1 FILLER_0_27_896 ();
 sg13g2_fill_2 FILLER_0_27_902 ();
 sg13g2_fill_2 FILLER_0_27_930 ();
 sg13g2_fill_1 FILLER_0_27_932 ();
 sg13g2_fill_2 FILLER_0_27_959 ();
 sg13g2_fill_4 FILLER_0_27_966 ();
 sg13g2_fill_2 FILLER_0_27_970 ();
 sg13g2_fill_8 FILLER_0_27_998 ();
 sg13g2_fill_2 FILLER_0_27_1006 ();
 sg13g2_fill_1 FILLER_0_27_1008 ();
 sg13g2_fill_8 FILLER_0_27_1014 ();
 sg13g2_fill_8 FILLER_0_27_1022 ();
 sg13g2_fill_8 FILLER_0_27_1030 ();
 sg13g2_fill_8 FILLER_0_27_1038 ();
 sg13g2_fill_2 FILLER_0_27_1046 ();
 sg13g2_fill_2 FILLER_0_27_1053 ();
 sg13g2_fill_4 FILLER_0_27_1062 ();
 sg13g2_fill_2 FILLER_0_27_1071 ();
 sg13g2_fill_8 FILLER_0_27_1099 ();
 sg13g2_fill_8 FILLER_0_27_1107 ();
 sg13g2_fill_8 FILLER_0_27_1115 ();
 sg13g2_fill_8 FILLER_0_27_1123 ();
 sg13g2_fill_8 FILLER_0_27_1131 ();
 sg13g2_fill_8 FILLER_0_27_1139 ();
 sg13g2_fill_2 FILLER_0_27_1147 ();
 sg13g2_fill_2 FILLER_0_27_1157 ();
 sg13g2_fill_2 FILLER_0_27_1164 ();
 sg13g2_fill_2 FILLER_0_27_1173 ();
 sg13g2_fill_4 FILLER_0_27_1179 ();
 sg13g2_fill_2 FILLER_0_27_1183 ();
 sg13g2_fill_2 FILLER_0_27_1192 ();
 sg13g2_fill_2 FILLER_0_27_1199 ();
 sg13g2_fill_4 FILLER_0_27_1209 ();
 sg13g2_fill_1 FILLER_0_27_1213 ();
 sg13g2_fill_2 FILLER_0_27_1222 ();
 sg13g2_fill_8 FILLER_0_27_1229 ();
 sg13g2_fill_8 FILLER_0_27_1237 ();
 sg13g2_fill_4 FILLER_0_27_1245 ();
 sg13g2_fill_8 FILLER_0_27_1259 ();
 sg13g2_fill_8 FILLER_0_27_1267 ();
 sg13g2_fill_4 FILLER_0_27_1275 ();
 sg13g2_fill_8 FILLER_0_27_1287 ();
 sg13g2_fill_2 FILLER_0_27_1295 ();
 sg13g2_fill_8 FILLER_0_28_0 ();
 sg13g2_fill_8 FILLER_0_28_8 ();
 sg13g2_fill_8 FILLER_0_28_16 ();
 sg13g2_fill_8 FILLER_0_28_24 ();
 sg13g2_fill_8 FILLER_0_28_32 ();
 sg13g2_fill_8 FILLER_0_28_40 ();
 sg13g2_fill_8 FILLER_0_28_48 ();
 sg13g2_fill_8 FILLER_0_28_56 ();
 sg13g2_fill_8 FILLER_0_28_64 ();
 sg13g2_fill_8 FILLER_0_28_72 ();
 sg13g2_fill_8 FILLER_0_28_80 ();
 sg13g2_fill_8 FILLER_0_28_88 ();
 sg13g2_fill_8 FILLER_0_28_96 ();
 sg13g2_fill_8 FILLER_0_28_104 ();
 sg13g2_fill_8 FILLER_0_28_112 ();
 sg13g2_fill_8 FILLER_0_28_120 ();
 sg13g2_fill_8 FILLER_0_28_128 ();
 sg13g2_fill_8 FILLER_0_28_136 ();
 sg13g2_fill_8 FILLER_0_28_144 ();
 sg13g2_fill_8 FILLER_0_28_152 ();
 sg13g2_fill_8 FILLER_0_28_160 ();
 sg13g2_fill_8 FILLER_0_28_168 ();
 sg13g2_fill_8 FILLER_0_28_176 ();
 sg13g2_fill_8 FILLER_0_28_184 ();
 sg13g2_fill_8 FILLER_0_28_192 ();
 sg13g2_fill_8 FILLER_0_28_200 ();
 sg13g2_fill_8 FILLER_0_28_208 ();
 sg13g2_fill_8 FILLER_0_28_216 ();
 sg13g2_fill_4 FILLER_0_28_224 ();
 sg13g2_fill_2 FILLER_0_28_228 ();
 sg13g2_fill_1 FILLER_0_28_230 ();
 sg13g2_fill_2 FILLER_0_28_236 ();
 sg13g2_fill_1 FILLER_0_28_238 ();
 sg13g2_fill_4 FILLER_0_28_243 ();
 sg13g2_fill_2 FILLER_0_28_247 ();
 sg13g2_fill_1 FILLER_0_28_249 ();
 sg13g2_fill_4 FILLER_0_28_271 ();
 sg13g2_fill_2 FILLER_0_28_275 ();
 sg13g2_fill_8 FILLER_0_28_282 ();
 sg13g2_fill_4 FILLER_0_28_290 ();
 sg13g2_fill_2 FILLER_0_28_294 ();
 sg13g2_fill_1 FILLER_0_28_296 ();
 sg13g2_fill_2 FILLER_0_28_301 ();
 sg13g2_fill_4 FILLER_0_28_308 ();
 sg13g2_fill_2 FILLER_0_28_333 ();
 sg13g2_fill_2 FILLER_0_28_361 ();
 sg13g2_fill_8 FILLER_0_28_367 ();
 sg13g2_fill_4 FILLER_0_28_375 ();
 sg13g2_fill_1 FILLER_0_28_379 ();
 sg13g2_fill_8 FILLER_0_28_383 ();
 sg13g2_fill_8 FILLER_0_28_391 ();
 sg13g2_fill_8 FILLER_0_28_399 ();
 sg13g2_fill_4 FILLER_0_28_407 ();
 sg13g2_fill_2 FILLER_0_28_411 ();
 sg13g2_fill_2 FILLER_0_28_439 ();
 sg13g2_fill_2 FILLER_0_28_445 ();
 sg13g2_fill_1 FILLER_0_28_447 ();
 sg13g2_fill_8 FILLER_0_28_453 ();
 sg13g2_fill_8 FILLER_0_28_461 ();
 sg13g2_fill_8 FILLER_0_28_469 ();
 sg13g2_fill_4 FILLER_0_28_477 ();
 sg13g2_fill_2 FILLER_0_28_481 ();
 sg13g2_fill_2 FILLER_0_28_509 ();
 sg13g2_fill_2 FILLER_0_28_515 ();
 sg13g2_fill_8 FILLER_0_28_538 ();
 sg13g2_fill_4 FILLER_0_28_546 ();
 sg13g2_fill_2 FILLER_0_28_550 ();
 sg13g2_fill_1 FILLER_0_28_552 ();
 sg13g2_fill_2 FILLER_0_28_557 ();
 sg13g2_fill_2 FILLER_0_28_564 ();
 sg13g2_fill_2 FILLER_0_28_592 ();
 sg13g2_fill_8 FILLER_0_28_600 ();
 sg13g2_fill_8 FILLER_0_28_608 ();
 sg13g2_fill_8 FILLER_0_28_616 ();
 sg13g2_fill_8 FILLER_0_28_624 ();
 sg13g2_fill_4 FILLER_0_28_632 ();
 sg13g2_fill_8 FILLER_0_28_641 ();
 sg13g2_fill_8 FILLER_0_28_649 ();
 sg13g2_fill_8 FILLER_0_28_657 ();
 sg13g2_fill_4 FILLER_0_28_665 ();
 sg13g2_fill_2 FILLER_0_28_674 ();
 sg13g2_fill_2 FILLER_0_28_680 ();
 sg13g2_fill_2 FILLER_0_28_708 ();
 sg13g2_fill_2 FILLER_0_28_736 ();
 sg13g2_fill_2 FILLER_0_28_764 ();
 sg13g2_fill_2 FILLER_0_28_787 ();
 sg13g2_fill_2 FILLER_0_28_810 ();
 sg13g2_fill_8 FILLER_0_28_816 ();
 sg13g2_fill_2 FILLER_0_28_824 ();
 sg13g2_fill_1 FILLER_0_28_826 ();
 sg13g2_fill_8 FILLER_0_28_853 ();
 sg13g2_fill_8 FILLER_0_28_861 ();
 sg13g2_fill_1 FILLER_0_28_869 ();
 sg13g2_fill_8 FILLER_0_28_882 ();
 sg13g2_fill_1 FILLER_0_28_890 ();
 sg13g2_fill_4 FILLER_0_28_896 ();
 sg13g2_fill_8 FILLER_0_28_904 ();
 sg13g2_fill_4 FILLER_0_28_912 ();
 sg13g2_fill_2 FILLER_0_28_921 ();
 sg13g2_fill_8 FILLER_0_28_944 ();
 sg13g2_fill_1 FILLER_0_28_952 ();
 sg13g2_fill_2 FILLER_0_28_957 ();
 sg13g2_fill_2 FILLER_0_28_964 ();
 sg13g2_fill_1 FILLER_0_28_966 ();
 sg13g2_fill_4 FILLER_0_28_972 ();
 sg13g2_fill_8 FILLER_0_28_980 ();
 sg13g2_fill_1 FILLER_0_28_988 ();
 sg13g2_fill_8 FILLER_0_28_994 ();
 sg13g2_fill_8 FILLER_0_28_1002 ();
 sg13g2_fill_8 FILLER_0_28_1010 ();
 sg13g2_fill_8 FILLER_0_28_1018 ();
 sg13g2_fill_8 FILLER_0_28_1026 ();
 sg13g2_fill_8 FILLER_0_28_1034 ();
 sg13g2_fill_4 FILLER_0_28_1042 ();
 sg13g2_fill_2 FILLER_0_28_1046 ();
 sg13g2_fill_1 FILLER_0_28_1048 ();
 sg13g2_fill_8 FILLER_0_28_1057 ();
 sg13g2_fill_4 FILLER_0_28_1065 ();
 sg13g2_fill_1 FILLER_0_28_1069 ();
 sg13g2_fill_4 FILLER_0_28_1074 ();
 sg13g2_fill_1 FILLER_0_28_1078 ();
 sg13g2_fill_4 FILLER_0_28_1087 ();
 sg13g2_fill_1 FILLER_0_28_1091 ();
 sg13g2_fill_8 FILLER_0_28_1113 ();
 sg13g2_fill_8 FILLER_0_28_1121 ();
 sg13g2_fill_2 FILLER_0_28_1129 ();
 sg13g2_fill_1 FILLER_0_28_1131 ();
 sg13g2_fill_8 FILLER_0_28_1136 ();
 sg13g2_fill_4 FILLER_0_28_1144 ();
 sg13g2_fill_2 FILLER_0_28_1148 ();
 sg13g2_fill_1 FILLER_0_28_1150 ();
 sg13g2_fill_2 FILLER_0_28_1155 ();
 sg13g2_fill_2 FILLER_0_28_1165 ();
 sg13g2_fill_1 FILLER_0_28_1167 ();
 sg13g2_fill_2 FILLER_0_28_1174 ();
 sg13g2_fill_1 FILLER_0_28_1176 ();
 sg13g2_fill_4 FILLER_0_28_1182 ();
 sg13g2_fill_1 FILLER_0_28_1186 ();
 sg13g2_fill_2 FILLER_0_28_1192 ();
 sg13g2_fill_8 FILLER_0_28_1198 ();
 sg13g2_fill_2 FILLER_0_28_1206 ();
 sg13g2_fill_1 FILLER_0_28_1208 ();
 sg13g2_fill_2 FILLER_0_28_1214 ();
 sg13g2_fill_1 FILLER_0_28_1216 ();
 sg13g2_fill_2 FILLER_0_28_1221 ();
 sg13g2_fill_8 FILLER_0_28_1227 ();
 sg13g2_fill_8 FILLER_0_28_1235 ();
 sg13g2_fill_8 FILLER_0_28_1243 ();
 sg13g2_fill_4 FILLER_0_28_1251 ();
 sg13g2_fill_1 FILLER_0_28_1255 ();
 sg13g2_fill_8 FILLER_0_28_1261 ();
 sg13g2_fill_8 FILLER_0_28_1269 ();
 sg13g2_fill_2 FILLER_0_28_1277 ();
 sg13g2_fill_8 FILLER_0_28_1286 ();
 sg13g2_fill_2 FILLER_0_28_1294 ();
 sg13g2_fill_1 FILLER_0_28_1296 ();
 sg13g2_fill_8 FILLER_0_29_0 ();
 sg13g2_fill_8 FILLER_0_29_8 ();
 sg13g2_fill_8 FILLER_0_29_16 ();
 sg13g2_fill_8 FILLER_0_29_24 ();
 sg13g2_fill_8 FILLER_0_29_32 ();
 sg13g2_fill_8 FILLER_0_29_40 ();
 sg13g2_fill_8 FILLER_0_29_48 ();
 sg13g2_fill_8 FILLER_0_29_56 ();
 sg13g2_fill_8 FILLER_0_29_64 ();
 sg13g2_fill_8 FILLER_0_29_72 ();
 sg13g2_fill_8 FILLER_0_29_80 ();
 sg13g2_fill_8 FILLER_0_29_88 ();
 sg13g2_fill_8 FILLER_0_29_96 ();
 sg13g2_fill_8 FILLER_0_29_104 ();
 sg13g2_fill_8 FILLER_0_29_112 ();
 sg13g2_fill_8 FILLER_0_29_120 ();
 sg13g2_fill_8 FILLER_0_29_128 ();
 sg13g2_fill_8 FILLER_0_29_136 ();
 sg13g2_fill_8 FILLER_0_29_144 ();
 sg13g2_fill_8 FILLER_0_29_152 ();
 sg13g2_fill_8 FILLER_0_29_160 ();
 sg13g2_fill_8 FILLER_0_29_168 ();
 sg13g2_fill_8 FILLER_0_29_176 ();
 sg13g2_fill_8 FILLER_0_29_184 ();
 sg13g2_fill_8 FILLER_0_29_192 ();
 sg13g2_fill_8 FILLER_0_29_200 ();
 sg13g2_fill_8 FILLER_0_29_208 ();
 sg13g2_fill_8 FILLER_0_29_216 ();
 sg13g2_fill_8 FILLER_0_29_224 ();
 sg13g2_fill_8 FILLER_0_29_232 ();
 sg13g2_fill_8 FILLER_0_29_240 ();
 sg13g2_fill_8 FILLER_0_29_248 ();
 sg13g2_fill_8 FILLER_0_29_256 ();
 sg13g2_fill_8 FILLER_0_29_264 ();
 sg13g2_fill_8 FILLER_0_29_272 ();
 sg13g2_fill_8 FILLER_0_29_280 ();
 sg13g2_fill_8 FILLER_0_29_288 ();
 sg13g2_fill_8 FILLER_0_29_296 ();
 sg13g2_fill_8 FILLER_0_29_304 ();
 sg13g2_fill_8 FILLER_0_29_312 ();
 sg13g2_fill_8 FILLER_0_29_320 ();
 sg13g2_fill_8 FILLER_0_29_328 ();
 sg13g2_fill_8 FILLER_0_29_336 ();
 sg13g2_fill_8 FILLER_0_29_344 ();
 sg13g2_fill_8 FILLER_0_29_352 ();
 sg13g2_fill_8 FILLER_0_29_360 ();
 sg13g2_fill_8 FILLER_0_29_368 ();
 sg13g2_fill_8 FILLER_0_29_376 ();
 sg13g2_fill_8 FILLER_0_29_384 ();
 sg13g2_fill_8 FILLER_0_29_392 ();
 sg13g2_fill_2 FILLER_0_29_400 ();
 sg13g2_fill_8 FILLER_0_29_407 ();
 sg13g2_fill_1 FILLER_0_29_415 ();
 sg13g2_fill_2 FILLER_0_29_421 ();
 sg13g2_fill_8 FILLER_0_29_428 ();
 sg13g2_fill_8 FILLER_0_29_436 ();
 sg13g2_fill_8 FILLER_0_29_444 ();
 sg13g2_fill_8 FILLER_0_29_452 ();
 sg13g2_fill_8 FILLER_0_29_460 ();
 sg13g2_fill_8 FILLER_0_29_468 ();
 sg13g2_fill_8 FILLER_0_29_476 ();
 sg13g2_fill_2 FILLER_0_29_484 ();
 sg13g2_fill_4 FILLER_0_29_490 ();
 sg13g2_fill_1 FILLER_0_29_494 ();
 sg13g2_fill_8 FILLER_0_29_499 ();
 sg13g2_fill_1 FILLER_0_29_507 ();
 sg13g2_fill_2 FILLER_0_29_518 ();
 sg13g2_fill_8 FILLER_0_29_525 ();
 sg13g2_fill_8 FILLER_0_29_533 ();
 sg13g2_fill_2 FILLER_0_29_546 ();
 sg13g2_fill_2 FILLER_0_29_556 ();
 sg13g2_fill_8 FILLER_0_29_562 ();
 sg13g2_fill_8 FILLER_0_29_570 ();
 sg13g2_fill_8 FILLER_0_29_578 ();
 sg13g2_fill_8 FILLER_0_29_586 ();
 sg13g2_fill_8 FILLER_0_29_594 ();
 sg13g2_fill_2 FILLER_0_29_602 ();
 sg13g2_fill_1 FILLER_0_29_604 ();
 sg13g2_fill_8 FILLER_0_29_609 ();
 sg13g2_fill_8 FILLER_0_29_617 ();
 sg13g2_fill_4 FILLER_0_29_625 ();
 sg13g2_fill_2 FILLER_0_29_629 ();
 sg13g2_fill_1 FILLER_0_29_631 ();
 sg13g2_fill_4 FILLER_0_29_637 ();
 sg13g2_fill_2 FILLER_0_29_645 ();
 sg13g2_fill_2 FILLER_0_29_673 ();
 sg13g2_fill_2 FILLER_0_29_680 ();
 sg13g2_fill_2 FILLER_0_29_687 ();
 sg13g2_fill_2 FILLER_0_29_693 ();
 sg13g2_fill_8 FILLER_0_29_716 ();
 sg13g2_fill_4 FILLER_0_29_724 ();
 sg13g2_fill_8 FILLER_0_29_732 ();
 sg13g2_fill_4 FILLER_0_29_745 ();
 sg13g2_fill_2 FILLER_0_29_754 ();
 sg13g2_fill_8 FILLER_0_29_760 ();
 sg13g2_fill_8 FILLER_0_29_768 ();
 sg13g2_fill_8 FILLER_0_29_776 ();
 sg13g2_fill_8 FILLER_0_29_784 ();
 sg13g2_fill_8 FILLER_0_29_792 ();
 sg13g2_fill_2 FILLER_0_29_800 ();
 sg13g2_fill_1 FILLER_0_29_802 ();
 sg13g2_fill_2 FILLER_0_29_808 ();
 sg13g2_fill_8 FILLER_0_29_815 ();
 sg13g2_fill_8 FILLER_0_29_823 ();
 sg13g2_fill_1 FILLER_0_29_831 ();
 sg13g2_fill_2 FILLER_0_29_837 ();
 sg13g2_fill_4 FILLER_0_29_843 ();
 sg13g2_fill_2 FILLER_0_29_853 ();
 sg13g2_fill_8 FILLER_0_29_860 ();
 sg13g2_fill_8 FILLER_0_29_868 ();
 sg13g2_fill_4 FILLER_0_29_876 ();
 sg13g2_fill_2 FILLER_0_29_880 ();
 sg13g2_fill_8 FILLER_0_29_908 ();
 sg13g2_fill_8 FILLER_0_29_916 ();
 sg13g2_fill_8 FILLER_0_29_924 ();
 sg13g2_fill_8 FILLER_0_29_932 ();
 sg13g2_fill_8 FILLER_0_29_940 ();
 sg13g2_fill_8 FILLER_0_29_948 ();
 sg13g2_fill_2 FILLER_0_29_956 ();
 sg13g2_fill_4 FILLER_0_29_964 ();
 sg13g2_fill_2 FILLER_0_29_968 ();
 sg13g2_fill_8 FILLER_0_29_975 ();
 sg13g2_fill_8 FILLER_0_29_983 ();
 sg13g2_fill_8 FILLER_0_29_991 ();
 sg13g2_fill_1 FILLER_0_29_999 ();
 sg13g2_fill_2 FILLER_0_29_1004 ();
 sg13g2_fill_2 FILLER_0_29_1011 ();
 sg13g2_fill_8 FILLER_0_29_1039 ();
 sg13g2_fill_8 FILLER_0_29_1047 ();
 sg13g2_fill_8 FILLER_0_29_1055 ();
 sg13g2_fill_8 FILLER_0_29_1063 ();
 sg13g2_fill_4 FILLER_0_29_1071 ();
 sg13g2_fill_2 FILLER_0_29_1075 ();
 sg13g2_fill_1 FILLER_0_29_1077 ();
 sg13g2_fill_2 FILLER_0_29_1083 ();
 sg13g2_fill_4 FILLER_0_29_1090 ();
 sg13g2_fill_2 FILLER_0_29_1094 ();
 sg13g2_fill_1 FILLER_0_29_1096 ();
 sg13g2_fill_2 FILLER_0_29_1101 ();
 sg13g2_fill_4 FILLER_0_29_1129 ();
 sg13g2_fill_2 FILLER_0_29_1133 ();
 sg13g2_fill_4 FILLER_0_29_1139 ();
 sg13g2_fill_2 FILLER_0_29_1151 ();
 sg13g2_fill_8 FILLER_0_29_1158 ();
 sg13g2_fill_2 FILLER_0_29_1171 ();
 sg13g2_fill_8 FILLER_0_29_1178 ();
 sg13g2_fill_8 FILLER_0_29_1186 ();
 sg13g2_fill_8 FILLER_0_29_1194 ();
 sg13g2_fill_8 FILLER_0_29_1202 ();
 sg13g2_fill_8 FILLER_0_29_1210 ();
 sg13g2_fill_8 FILLER_0_29_1218 ();
 sg13g2_fill_8 FILLER_0_29_1226 ();
 sg13g2_fill_8 FILLER_0_29_1234 ();
 sg13g2_fill_4 FILLER_0_29_1242 ();
 sg13g2_fill_2 FILLER_0_29_1246 ();
 sg13g2_fill_1 FILLER_0_29_1248 ();
 sg13g2_fill_4 FILLER_0_29_1254 ();
 sg13g2_fill_2 FILLER_0_29_1258 ();
 sg13g2_fill_1 FILLER_0_29_1260 ();
 sg13g2_fill_8 FILLER_0_29_1269 ();
 sg13g2_fill_1 FILLER_0_29_1277 ();
 sg13g2_fill_2 FILLER_0_29_1283 ();
 sg13g2_fill_8 FILLER_0_29_1289 ();
 sg13g2_fill_8 FILLER_0_30_0 ();
 sg13g2_fill_8 FILLER_0_30_8 ();
 sg13g2_fill_8 FILLER_0_30_16 ();
 sg13g2_fill_8 FILLER_0_30_24 ();
 sg13g2_fill_8 FILLER_0_30_32 ();
 sg13g2_fill_8 FILLER_0_30_40 ();
 sg13g2_fill_8 FILLER_0_30_48 ();
 sg13g2_fill_8 FILLER_0_30_56 ();
 sg13g2_fill_8 FILLER_0_30_64 ();
 sg13g2_fill_8 FILLER_0_30_72 ();
 sg13g2_fill_8 FILLER_0_30_80 ();
 sg13g2_fill_8 FILLER_0_30_88 ();
 sg13g2_fill_8 FILLER_0_30_96 ();
 sg13g2_fill_8 FILLER_0_30_104 ();
 sg13g2_fill_8 FILLER_0_30_112 ();
 sg13g2_fill_8 FILLER_0_30_120 ();
 sg13g2_fill_8 FILLER_0_30_128 ();
 sg13g2_fill_8 FILLER_0_30_136 ();
 sg13g2_fill_8 FILLER_0_30_144 ();
 sg13g2_fill_8 FILLER_0_30_152 ();
 sg13g2_fill_8 FILLER_0_30_160 ();
 sg13g2_fill_8 FILLER_0_30_168 ();
 sg13g2_fill_8 FILLER_0_30_176 ();
 sg13g2_fill_8 FILLER_0_30_184 ();
 sg13g2_fill_8 FILLER_0_30_192 ();
 sg13g2_fill_4 FILLER_0_30_200 ();
 sg13g2_fill_1 FILLER_0_30_204 ();
 sg13g2_fill_2 FILLER_0_30_231 ();
 sg13g2_fill_2 FILLER_0_30_238 ();
 sg13g2_fill_1 FILLER_0_30_240 ();
 sg13g2_fill_8 FILLER_0_30_245 ();
 sg13g2_fill_8 FILLER_0_30_253 ();
 sg13g2_fill_8 FILLER_0_30_261 ();
 sg13g2_fill_8 FILLER_0_30_269 ();
 sg13g2_fill_8 FILLER_0_30_277 ();
 sg13g2_fill_2 FILLER_0_30_285 ();
 sg13g2_fill_1 FILLER_0_30_287 ();
 sg13g2_fill_2 FILLER_0_30_293 ();
 sg13g2_fill_8 FILLER_0_30_299 ();
 sg13g2_fill_8 FILLER_0_30_307 ();
 sg13g2_fill_8 FILLER_0_30_315 ();
 sg13g2_fill_8 FILLER_0_30_323 ();
 sg13g2_fill_8 FILLER_0_30_331 ();
 sg13g2_fill_8 FILLER_0_30_339 ();
 sg13g2_fill_8 FILLER_0_30_347 ();
 sg13g2_fill_4 FILLER_0_30_355 ();
 sg13g2_fill_2 FILLER_0_30_363 ();
 sg13g2_fill_8 FILLER_0_30_371 ();
 sg13g2_fill_1 FILLER_0_30_379 ();
 sg13g2_fill_8 FILLER_0_30_385 ();
 sg13g2_fill_4 FILLER_0_30_393 ();
 sg13g2_fill_1 FILLER_0_30_397 ();
 sg13g2_fill_8 FILLER_0_30_403 ();
 sg13g2_fill_8 FILLER_0_30_411 ();
 sg13g2_fill_8 FILLER_0_30_419 ();
 sg13g2_fill_8 FILLER_0_30_427 ();
 sg13g2_fill_8 FILLER_0_30_435 ();
 sg13g2_fill_4 FILLER_0_30_443 ();
 sg13g2_fill_8 FILLER_0_30_452 ();
 sg13g2_fill_8 FILLER_0_30_460 ();
 sg13g2_fill_8 FILLER_0_30_468 ();
 sg13g2_fill_8 FILLER_0_30_476 ();
 sg13g2_fill_4 FILLER_0_30_484 ();
 sg13g2_fill_1 FILLER_0_30_488 ();
 sg13g2_fill_8 FILLER_0_30_494 ();
 sg13g2_fill_4 FILLER_0_30_502 ();
 sg13g2_fill_1 FILLER_0_30_506 ();
 sg13g2_fill_4 FILLER_0_30_512 ();
 sg13g2_fill_2 FILLER_0_30_516 ();
 sg13g2_fill_2 FILLER_0_30_523 ();
 sg13g2_fill_2 FILLER_0_30_529 ();
 sg13g2_fill_4 FILLER_0_30_541 ();
 sg13g2_fill_4 FILLER_0_30_550 ();
 sg13g2_fill_2 FILLER_0_30_554 ();
 sg13g2_fill_1 FILLER_0_30_556 ();
 sg13g2_fill_8 FILLER_0_30_561 ();
 sg13g2_fill_8 FILLER_0_30_569 ();
 sg13g2_fill_8 FILLER_0_30_577 ();
 sg13g2_fill_8 FILLER_0_30_585 ();
 sg13g2_fill_4 FILLER_0_30_593 ();
 sg13g2_fill_2 FILLER_0_30_597 ();
 sg13g2_fill_2 FILLER_0_30_604 ();
 sg13g2_fill_8 FILLER_0_30_610 ();
 sg13g2_fill_8 FILLER_0_30_618 ();
 sg13g2_fill_8 FILLER_0_30_626 ();
 sg13g2_fill_8 FILLER_0_30_634 ();
 sg13g2_fill_8 FILLER_0_30_642 ();
 sg13g2_fill_8 FILLER_0_30_650 ();
 sg13g2_fill_8 FILLER_0_30_658 ();
 sg13g2_fill_8 FILLER_0_30_666 ();
 sg13g2_fill_8 FILLER_0_30_674 ();
 sg13g2_fill_1 FILLER_0_30_682 ();
 sg13g2_fill_8 FILLER_0_30_691 ();
 sg13g2_fill_4 FILLER_0_30_699 ();
 sg13g2_fill_2 FILLER_0_30_703 ();
 sg13g2_fill_1 FILLER_0_30_705 ();
 sg13g2_fill_8 FILLER_0_30_711 ();
 sg13g2_fill_8 FILLER_0_30_719 ();
 sg13g2_fill_8 FILLER_0_30_727 ();
 sg13g2_fill_8 FILLER_0_30_735 ();
 sg13g2_fill_8 FILLER_0_30_743 ();
 sg13g2_fill_8 FILLER_0_30_751 ();
 sg13g2_fill_8 FILLER_0_30_759 ();
 sg13g2_fill_8 FILLER_0_30_767 ();
 sg13g2_fill_8 FILLER_0_30_775 ();
 sg13g2_fill_8 FILLER_0_30_783 ();
 sg13g2_fill_8 FILLER_0_30_795 ();
 sg13g2_fill_8 FILLER_0_30_803 ();
 sg13g2_fill_8 FILLER_0_30_811 ();
 sg13g2_fill_8 FILLER_0_30_819 ();
 sg13g2_fill_8 FILLER_0_30_827 ();
 sg13g2_fill_8 FILLER_0_30_835 ();
 sg13g2_fill_8 FILLER_0_30_843 ();
 sg13g2_fill_8 FILLER_0_30_851 ();
 sg13g2_fill_4 FILLER_0_30_859 ();
 sg13g2_fill_1 FILLER_0_30_863 ();
 sg13g2_fill_2 FILLER_0_30_869 ();
 sg13g2_fill_8 FILLER_0_30_875 ();
 sg13g2_fill_8 FILLER_0_30_883 ();
 sg13g2_fill_8 FILLER_0_30_912 ();
 sg13g2_fill_8 FILLER_0_30_920 ();
 sg13g2_fill_4 FILLER_0_30_928 ();
 sg13g2_fill_1 FILLER_0_30_932 ();
 sg13g2_fill_8 FILLER_0_30_938 ();
 sg13g2_fill_2 FILLER_0_30_972 ();
 sg13g2_fill_8 FILLER_0_30_984 ();
 sg13g2_fill_8 FILLER_0_30_992 ();
 sg13g2_fill_8 FILLER_0_30_1000 ();
 sg13g2_fill_8 FILLER_0_30_1008 ();
 sg13g2_fill_1 FILLER_0_30_1016 ();
 sg13g2_fill_2 FILLER_0_30_1024 ();
 sg13g2_fill_8 FILLER_0_30_1047 ();
 sg13g2_fill_8 FILLER_0_30_1055 ();
 sg13g2_fill_8 FILLER_0_30_1063 ();
 sg13g2_fill_8 FILLER_0_30_1071 ();
 sg13g2_fill_4 FILLER_0_30_1079 ();
 sg13g2_fill_1 FILLER_0_30_1083 ();
 sg13g2_fill_2 FILLER_0_30_1088 ();
 sg13g2_fill_8 FILLER_0_30_1111 ();
 sg13g2_fill_1 FILLER_0_30_1119 ();
 sg13g2_fill_2 FILLER_0_30_1125 ();
 sg13g2_fill_4 FILLER_0_30_1132 ();
 sg13g2_fill_1 FILLER_0_30_1136 ();
 sg13g2_fill_2 FILLER_0_30_1142 ();
 sg13g2_fill_4 FILLER_0_30_1148 ();
 sg13g2_fill_8 FILLER_0_30_1158 ();
 sg13g2_fill_8 FILLER_0_30_1166 ();
 sg13g2_fill_8 FILLER_0_30_1174 ();
 sg13g2_fill_8 FILLER_0_30_1182 ();
 sg13g2_fill_8 FILLER_0_30_1190 ();
 sg13g2_fill_8 FILLER_0_30_1198 ();
 sg13g2_fill_8 FILLER_0_30_1206 ();
 sg13g2_fill_2 FILLER_0_30_1218 ();
 sg13g2_fill_1 FILLER_0_30_1220 ();
 sg13g2_fill_2 FILLER_0_30_1247 ();
 sg13g2_fill_2 FILLER_0_30_1254 ();
 sg13g2_fill_2 FILLER_0_30_1282 ();
 sg13g2_fill_8 FILLER_0_30_1288 ();
 sg13g2_fill_1 FILLER_0_30_1296 ();
 sg13g2_fill_8 FILLER_0_31_0 ();
 sg13g2_fill_8 FILLER_0_31_8 ();
 sg13g2_fill_8 FILLER_0_31_16 ();
 sg13g2_fill_8 FILLER_0_31_24 ();
 sg13g2_fill_8 FILLER_0_31_32 ();
 sg13g2_fill_8 FILLER_0_31_40 ();
 sg13g2_fill_8 FILLER_0_31_48 ();
 sg13g2_fill_8 FILLER_0_31_56 ();
 sg13g2_fill_8 FILLER_0_31_64 ();
 sg13g2_fill_8 FILLER_0_31_72 ();
 sg13g2_fill_8 FILLER_0_31_80 ();
 sg13g2_fill_8 FILLER_0_31_88 ();
 sg13g2_fill_8 FILLER_0_31_96 ();
 sg13g2_fill_8 FILLER_0_31_104 ();
 sg13g2_fill_8 FILLER_0_31_112 ();
 sg13g2_fill_8 FILLER_0_31_120 ();
 sg13g2_fill_8 FILLER_0_31_128 ();
 sg13g2_fill_8 FILLER_0_31_136 ();
 sg13g2_fill_8 FILLER_0_31_144 ();
 sg13g2_fill_8 FILLER_0_31_152 ();
 sg13g2_fill_8 FILLER_0_31_160 ();
 sg13g2_fill_8 FILLER_0_31_168 ();
 sg13g2_fill_8 FILLER_0_31_176 ();
 sg13g2_fill_8 FILLER_0_31_184 ();
 sg13g2_fill_8 FILLER_0_31_192 ();
 sg13g2_fill_8 FILLER_0_31_200 ();
 sg13g2_fill_2 FILLER_0_31_208 ();
 sg13g2_fill_1 FILLER_0_31_210 ();
 sg13g2_fill_2 FILLER_0_31_216 ();
 sg13g2_fill_2 FILLER_0_31_222 ();
 sg13g2_fill_1 FILLER_0_31_224 ();
 sg13g2_fill_8 FILLER_0_31_251 ();
 sg13g2_fill_4 FILLER_0_31_259 ();
 sg13g2_fill_2 FILLER_0_31_267 ();
 sg13g2_fill_2 FILLER_0_31_274 ();
 sg13g2_fill_4 FILLER_0_31_280 ();
 sg13g2_fill_2 FILLER_0_31_284 ();
 sg13g2_fill_1 FILLER_0_31_286 ();
 sg13g2_fill_8 FILLER_0_31_313 ();
 sg13g2_fill_8 FILLER_0_31_321 ();
 sg13g2_fill_8 FILLER_0_31_329 ();
 sg13g2_fill_4 FILLER_0_31_337 ();
 sg13g2_fill_1 FILLER_0_31_341 ();
 sg13g2_fill_2 FILLER_0_31_368 ();
 sg13g2_fill_8 FILLER_0_31_378 ();
 sg13g2_fill_4 FILLER_0_31_390 ();
 sg13g2_fill_1 FILLER_0_31_394 ();
 sg13g2_fill_8 FILLER_0_31_402 ();
 sg13g2_fill_8 FILLER_0_31_410 ();
 sg13g2_fill_8 FILLER_0_31_418 ();
 sg13g2_fill_8 FILLER_0_31_426 ();
 sg13g2_fill_8 FILLER_0_31_434 ();
 sg13g2_fill_4 FILLER_0_31_442 ();
 sg13g2_fill_2 FILLER_0_31_446 ();
 sg13g2_fill_2 FILLER_0_31_453 ();
 sg13g2_fill_8 FILLER_0_31_476 ();
 sg13g2_fill_8 FILLER_0_31_484 ();
 sg13g2_fill_4 FILLER_0_31_492 ();
 sg13g2_fill_4 FILLER_0_31_500 ();
 sg13g2_fill_8 FILLER_0_31_530 ();
 sg13g2_fill_8 FILLER_0_31_538 ();
 sg13g2_fill_4 FILLER_0_31_546 ();
 sg13g2_fill_2 FILLER_0_31_550 ();
 sg13g2_fill_1 FILLER_0_31_552 ();
 sg13g2_fill_8 FILLER_0_31_557 ();
 sg13g2_fill_8 FILLER_0_31_565 ();
 sg13g2_fill_8 FILLER_0_31_573 ();
 sg13g2_fill_8 FILLER_0_31_581 ();
 sg13g2_fill_8 FILLER_0_31_589 ();
 sg13g2_fill_4 FILLER_0_31_597 ();
 sg13g2_fill_2 FILLER_0_31_601 ();
 sg13g2_fill_1 FILLER_0_31_603 ();
 sg13g2_fill_2 FILLER_0_31_609 ();
 sg13g2_fill_8 FILLER_0_31_621 ();
 sg13g2_fill_8 FILLER_0_31_629 ();
 sg13g2_fill_8 FILLER_0_31_637 ();
 sg13g2_fill_2 FILLER_0_31_645 ();
 sg13g2_fill_1 FILLER_0_31_647 ();
 sg13g2_fill_2 FILLER_0_31_653 ();
 sg13g2_fill_8 FILLER_0_31_659 ();
 sg13g2_fill_8 FILLER_0_31_667 ();
 sg13g2_fill_8 FILLER_0_31_675 ();
 sg13g2_fill_8 FILLER_0_31_683 ();
 sg13g2_fill_8 FILLER_0_31_691 ();
 sg13g2_fill_8 FILLER_0_31_699 ();
 sg13g2_fill_8 FILLER_0_31_707 ();
 sg13g2_fill_8 FILLER_0_31_715 ();
 sg13g2_fill_8 FILLER_0_31_723 ();
 sg13g2_fill_4 FILLER_0_31_731 ();
 sg13g2_fill_8 FILLER_0_31_740 ();
 sg13g2_fill_8 FILLER_0_31_748 ();
 sg13g2_fill_8 FILLER_0_31_756 ();
 sg13g2_fill_8 FILLER_0_31_764 ();
 sg13g2_fill_2 FILLER_0_31_772 ();
 sg13g2_fill_1 FILLER_0_31_774 ();
 sg13g2_fill_2 FILLER_0_31_780 ();
 sg13g2_fill_2 FILLER_0_31_808 ();
 sg13g2_fill_8 FILLER_0_31_814 ();
 sg13g2_fill_8 FILLER_0_31_822 ();
 sg13g2_fill_8 FILLER_0_31_830 ();
 sg13g2_fill_8 FILLER_0_31_838 ();
 sg13g2_fill_8 FILLER_0_31_846 ();
 sg13g2_fill_4 FILLER_0_31_854 ();
 sg13g2_fill_2 FILLER_0_31_858 ();
 sg13g2_fill_1 FILLER_0_31_860 ();
 sg13g2_fill_2 FILLER_0_31_887 ();
 sg13g2_fill_2 FILLER_0_31_910 ();
 sg13g2_fill_8 FILLER_0_31_919 ();
 sg13g2_fill_8 FILLER_0_31_927 ();
 sg13g2_fill_8 FILLER_0_31_935 ();
 sg13g2_fill_4 FILLER_0_31_943 ();
 sg13g2_fill_2 FILLER_0_31_947 ();
 sg13g2_fill_1 FILLER_0_31_949 ();
 sg13g2_fill_2 FILLER_0_31_955 ();
 sg13g2_fill_8 FILLER_0_31_961 ();
 sg13g2_fill_8 FILLER_0_31_969 ();
 sg13g2_fill_4 FILLER_0_31_977 ();
 sg13g2_fill_1 FILLER_0_31_981 ();
 sg13g2_fill_2 FILLER_0_31_987 ();
 sg13g2_fill_8 FILLER_0_31_994 ();
 sg13g2_fill_2 FILLER_0_31_1007 ();
 sg13g2_fill_4 FILLER_0_31_1035 ();
 sg13g2_fill_8 FILLER_0_31_1044 ();
 sg13g2_fill_8 FILLER_0_31_1056 ();
 sg13g2_fill_2 FILLER_0_31_1090 ();
 sg13g2_fill_4 FILLER_0_31_1095 ();
 sg13g2_fill_8 FILLER_0_31_1104 ();
 sg13g2_fill_8 FILLER_0_31_1112 ();
 sg13g2_fill_8 FILLER_0_31_1120 ();
 sg13g2_fill_8 FILLER_0_31_1128 ();
 sg13g2_fill_8 FILLER_0_31_1136 ();
 sg13g2_fill_8 FILLER_0_31_1144 ();
 sg13g2_fill_8 FILLER_0_31_1152 ();
 sg13g2_fill_8 FILLER_0_31_1160 ();
 sg13g2_fill_8 FILLER_0_31_1168 ();
 sg13g2_fill_8 FILLER_0_31_1176 ();
 sg13g2_fill_8 FILLER_0_31_1184 ();
 sg13g2_fill_8 FILLER_0_31_1192 ();
 sg13g2_fill_8 FILLER_0_31_1200 ();
 sg13g2_fill_2 FILLER_0_31_1218 ();
 sg13g2_fill_8 FILLER_0_31_1225 ();
 sg13g2_fill_2 FILLER_0_31_1233 ();
 sg13g2_fill_1 FILLER_0_31_1235 ();
 sg13g2_fill_2 FILLER_0_31_1240 ();
 sg13g2_fill_2 FILLER_0_31_1247 ();
 sg13g2_fill_2 FILLER_0_31_1259 ();
 sg13g2_fill_2 FILLER_0_31_1266 ();
 sg13g2_fill_4 FILLER_0_31_1273 ();
 sg13g2_fill_2 FILLER_0_31_1277 ();
 sg13g2_fill_8 FILLER_0_31_1287 ();
 sg13g2_fill_2 FILLER_0_31_1295 ();
 sg13g2_fill_8 FILLER_0_32_0 ();
 sg13g2_fill_8 FILLER_0_32_8 ();
 sg13g2_fill_8 FILLER_0_32_16 ();
 sg13g2_fill_8 FILLER_0_32_24 ();
 sg13g2_fill_8 FILLER_0_32_32 ();
 sg13g2_fill_8 FILLER_0_32_40 ();
 sg13g2_fill_8 FILLER_0_32_48 ();
 sg13g2_fill_8 FILLER_0_32_56 ();
 sg13g2_fill_8 FILLER_0_32_64 ();
 sg13g2_fill_8 FILLER_0_32_72 ();
 sg13g2_fill_8 FILLER_0_32_80 ();
 sg13g2_fill_8 FILLER_0_32_88 ();
 sg13g2_fill_8 FILLER_0_32_96 ();
 sg13g2_fill_8 FILLER_0_32_104 ();
 sg13g2_fill_8 FILLER_0_32_112 ();
 sg13g2_fill_8 FILLER_0_32_120 ();
 sg13g2_fill_8 FILLER_0_32_128 ();
 sg13g2_fill_8 FILLER_0_32_136 ();
 sg13g2_fill_8 FILLER_0_32_144 ();
 sg13g2_fill_8 FILLER_0_32_152 ();
 sg13g2_fill_8 FILLER_0_32_160 ();
 sg13g2_fill_8 FILLER_0_32_168 ();
 sg13g2_fill_8 FILLER_0_32_176 ();
 sg13g2_fill_8 FILLER_0_32_184 ();
 sg13g2_fill_8 FILLER_0_32_192 ();
 sg13g2_fill_8 FILLER_0_32_200 ();
 sg13g2_fill_8 FILLER_0_32_208 ();
 sg13g2_fill_8 FILLER_0_32_216 ();
 sg13g2_fill_8 FILLER_0_32_224 ();
 sg13g2_fill_2 FILLER_0_32_232 ();
 sg13g2_fill_8 FILLER_0_32_255 ();
 sg13g2_fill_4 FILLER_0_32_263 ();
 sg13g2_fill_2 FILLER_0_32_267 ();
 sg13g2_fill_4 FILLER_0_32_295 ();
 sg13g2_fill_2 FILLER_0_32_299 ();
 sg13g2_fill_8 FILLER_0_32_322 ();
 sg13g2_fill_4 FILLER_0_32_330 ();
 sg13g2_fill_2 FILLER_0_32_339 ();
 sg13g2_fill_2 FILLER_0_32_346 ();
 sg13g2_fill_4 FILLER_0_32_352 ();
 sg13g2_fill_2 FILLER_0_32_360 ();
 sg13g2_fill_4 FILLER_0_32_367 ();
 sg13g2_fill_4 FILLER_0_32_376 ();
 sg13g2_fill_2 FILLER_0_32_380 ();
 sg13g2_fill_1 FILLER_0_32_382 ();
 sg13g2_fill_4 FILLER_0_32_388 ();
 sg13g2_fill_2 FILLER_0_32_392 ();
 sg13g2_fill_1 FILLER_0_32_394 ();
 sg13g2_fill_8 FILLER_0_32_400 ();
 sg13g2_fill_4 FILLER_0_32_408 ();
 sg13g2_fill_1 FILLER_0_32_412 ();
 sg13g2_fill_2 FILLER_0_32_418 ();
 sg13g2_fill_2 FILLER_0_32_425 ();
 sg13g2_fill_2 FILLER_0_32_431 ();
 sg13g2_fill_2 FILLER_0_32_437 ();
 sg13g2_fill_2 FILLER_0_32_465 ();
 sg13g2_fill_2 FILLER_0_32_472 ();
 sg13g2_fill_8 FILLER_0_32_478 ();
 sg13g2_fill_8 FILLER_0_32_486 ();
 sg13g2_fill_1 FILLER_0_32_494 ();
 sg13g2_fill_2 FILLER_0_32_500 ();
 sg13g2_fill_8 FILLER_0_32_528 ();
 sg13g2_fill_8 FILLER_0_32_536 ();
 sg13g2_fill_2 FILLER_0_32_544 ();
 sg13g2_fill_8 FILLER_0_32_551 ();
 sg13g2_fill_2 FILLER_0_32_559 ();
 sg13g2_fill_1 FILLER_0_32_561 ();
 sg13g2_fill_2 FILLER_0_32_566 ();
 sg13g2_fill_2 FILLER_0_32_573 ();
 sg13g2_fill_4 FILLER_0_32_601 ();
 sg13g2_fill_1 FILLER_0_32_605 ();
 sg13g2_fill_8 FILLER_0_32_632 ();
 sg13g2_fill_2 FILLER_0_32_666 ();
 sg13g2_fill_2 FILLER_0_32_673 ();
 sg13g2_fill_8 FILLER_0_32_679 ();
 sg13g2_fill_8 FILLER_0_32_687 ();
 sg13g2_fill_8 FILLER_0_32_695 ();
 sg13g2_fill_1 FILLER_0_32_703 ();
 sg13g2_fill_4 FILLER_0_32_708 ();
 sg13g2_fill_2 FILLER_0_32_712 ();
 sg13g2_fill_2 FILLER_0_32_719 ();
 sg13g2_fill_2 FILLER_0_32_725 ();
 sg13g2_fill_1 FILLER_0_32_727 ();
 sg13g2_fill_8 FILLER_0_32_732 ();
 sg13g2_fill_2 FILLER_0_32_740 ();
 sg13g2_fill_4 FILLER_0_32_746 ();
 sg13g2_fill_1 FILLER_0_32_750 ();
 sg13g2_fill_2 FILLER_0_32_756 ();
 sg13g2_fill_1 FILLER_0_32_758 ();
 sg13g2_fill_8 FILLER_0_32_763 ();
 sg13g2_fill_2 FILLER_0_32_771 ();
 sg13g2_fill_2 FILLER_0_32_799 ();
 sg13g2_fill_2 FILLER_0_32_806 ();
 sg13g2_fill_2 FILLER_0_32_813 ();
 sg13g2_fill_4 FILLER_0_32_819 ();
 sg13g2_fill_2 FILLER_0_32_823 ();
 sg13g2_fill_1 FILLER_0_32_825 ();
 sg13g2_fill_2 FILLER_0_32_831 ();
 sg13g2_fill_1 FILLER_0_32_833 ();
 sg13g2_fill_4 FILLER_0_32_855 ();
 sg13g2_fill_2 FILLER_0_32_859 ();
 sg13g2_fill_1 FILLER_0_32_861 ();
 sg13g2_fill_2 FILLER_0_32_888 ();
 sg13g2_fill_2 FILLER_0_32_894 ();
 sg13g2_fill_2 FILLER_0_32_922 ();
 sg13g2_fill_2 FILLER_0_32_929 ();
 sg13g2_fill_2 FILLER_0_32_937 ();
 sg13g2_fill_1 FILLER_0_32_939 ();
 sg13g2_fill_8 FILLER_0_32_945 ();
 sg13g2_fill_4 FILLER_0_32_953 ();
 sg13g2_fill_1 FILLER_0_32_957 ();
 sg13g2_fill_8 FILLER_0_32_963 ();
 sg13g2_fill_2 FILLER_0_32_971 ();
 sg13g2_fill_2 FILLER_0_32_978 ();
 sg13g2_fill_2 FILLER_0_32_985 ();
 sg13g2_fill_4 FILLER_0_32_994 ();
 sg13g2_fill_2 FILLER_0_32_998 ();
 sg13g2_fill_1 FILLER_0_32_1000 ();
 sg13g2_fill_2 FILLER_0_32_1005 ();
 sg13g2_fill_2 FILLER_0_32_1033 ();
 sg13g2_fill_4 FILLER_0_32_1061 ();
 sg13g2_fill_2 FILLER_0_32_1070 ();
 sg13g2_fill_8 FILLER_0_32_1076 ();
 sg13g2_fill_8 FILLER_0_32_1084 ();
 sg13g2_fill_8 FILLER_0_32_1092 ();
 sg13g2_fill_8 FILLER_0_32_1100 ();
 sg13g2_fill_8 FILLER_0_32_1108 ();
 sg13g2_fill_8 FILLER_0_32_1116 ();
 sg13g2_fill_4 FILLER_0_32_1124 ();
 sg13g2_fill_1 FILLER_0_32_1128 ();
 sg13g2_fill_2 FILLER_0_32_1137 ();
 sg13g2_fill_8 FILLER_0_32_1147 ();
 sg13g2_fill_8 FILLER_0_32_1155 ();
 sg13g2_fill_8 FILLER_0_32_1163 ();
 sg13g2_fill_8 FILLER_0_32_1171 ();
 sg13g2_fill_8 FILLER_0_32_1179 ();
 sg13g2_fill_8 FILLER_0_32_1187 ();
 sg13g2_fill_1 FILLER_0_32_1195 ();
 sg13g2_fill_4 FILLER_0_32_1200 ();
 sg13g2_fill_2 FILLER_0_32_1209 ();
 sg13g2_fill_8 FILLER_0_32_1215 ();
 sg13g2_fill_1 FILLER_0_32_1223 ();
 sg13g2_fill_8 FILLER_0_32_1229 ();
 sg13g2_fill_2 FILLER_0_32_1237 ();
 sg13g2_fill_1 FILLER_0_32_1239 ();
 sg13g2_fill_4 FILLER_0_32_1245 ();
 sg13g2_fill_2 FILLER_0_32_1249 ();
 sg13g2_fill_8 FILLER_0_32_1261 ();
 sg13g2_fill_8 FILLER_0_32_1269 ();
 sg13g2_fill_4 FILLER_0_32_1277 ();
 sg13g2_fill_8 FILLER_0_32_1285 ();
 sg13g2_fill_4 FILLER_0_32_1293 ();
 sg13g2_fill_8 FILLER_0_33_0 ();
 sg13g2_fill_8 FILLER_0_33_8 ();
 sg13g2_fill_8 FILLER_0_33_16 ();
 sg13g2_fill_8 FILLER_0_33_24 ();
 sg13g2_fill_8 FILLER_0_33_32 ();
 sg13g2_fill_8 FILLER_0_33_40 ();
 sg13g2_fill_8 FILLER_0_33_48 ();
 sg13g2_fill_8 FILLER_0_33_56 ();
 sg13g2_fill_8 FILLER_0_33_64 ();
 sg13g2_fill_8 FILLER_0_33_72 ();
 sg13g2_fill_8 FILLER_0_33_80 ();
 sg13g2_fill_8 FILLER_0_33_88 ();
 sg13g2_fill_8 FILLER_0_33_96 ();
 sg13g2_fill_8 FILLER_0_33_104 ();
 sg13g2_fill_8 FILLER_0_33_112 ();
 sg13g2_fill_8 FILLER_0_33_120 ();
 sg13g2_fill_8 FILLER_0_33_128 ();
 sg13g2_fill_8 FILLER_0_33_136 ();
 sg13g2_fill_8 FILLER_0_33_144 ();
 sg13g2_fill_8 FILLER_0_33_152 ();
 sg13g2_fill_8 FILLER_0_33_160 ();
 sg13g2_fill_8 FILLER_0_33_168 ();
 sg13g2_fill_8 FILLER_0_33_176 ();
 sg13g2_fill_8 FILLER_0_33_184 ();
 sg13g2_fill_8 FILLER_0_33_192 ();
 sg13g2_fill_8 FILLER_0_33_200 ();
 sg13g2_fill_4 FILLER_0_33_208 ();
 sg13g2_fill_8 FILLER_0_33_216 ();
 sg13g2_fill_8 FILLER_0_33_224 ();
 sg13g2_fill_1 FILLER_0_33_232 ();
 sg13g2_fill_4 FILLER_0_33_254 ();
 sg13g2_fill_2 FILLER_0_33_258 ();
 sg13g2_fill_2 FILLER_0_33_286 ();
 sg13g2_fill_8 FILLER_0_33_309 ();
 sg13g2_fill_8 FILLER_0_33_317 ();
 sg13g2_fill_8 FILLER_0_33_325 ();
 sg13g2_fill_4 FILLER_0_33_333 ();
 sg13g2_fill_2 FILLER_0_33_337 ();
 sg13g2_fill_2 FILLER_0_33_344 ();
 sg13g2_fill_8 FILLER_0_33_351 ();
 sg13g2_fill_8 FILLER_0_33_359 ();
 sg13g2_fill_8 FILLER_0_33_367 ();
 sg13g2_fill_4 FILLER_0_33_375 ();
 sg13g2_fill_1 FILLER_0_33_379 ();
 sg13g2_fill_8 FILLER_0_33_406 ();
 sg13g2_fill_4 FILLER_0_33_414 ();
 sg13g2_fill_1 FILLER_0_33_418 ();
 sg13g2_fill_4 FILLER_0_33_445 ();
 sg13g2_fill_1 FILLER_0_33_449 ();
 sg13g2_fill_2 FILLER_0_33_454 ();
 sg13g2_fill_1 FILLER_0_33_456 ();
 sg13g2_fill_8 FILLER_0_33_483 ();
 sg13g2_fill_8 FILLER_0_33_491 ();
 sg13g2_fill_8 FILLER_0_33_499 ();
 sg13g2_fill_8 FILLER_0_33_507 ();
 sg13g2_fill_8 FILLER_0_33_515 ();
 sg13g2_fill_8 FILLER_0_33_523 ();
 sg13g2_fill_8 FILLER_0_33_531 ();
 sg13g2_fill_4 FILLER_0_33_539 ();
 sg13g2_fill_1 FILLER_0_33_543 ();
 sg13g2_fill_2 FILLER_0_33_570 ();
 sg13g2_fill_1 FILLER_0_33_572 ();
 sg13g2_fill_8 FILLER_0_33_577 ();
 sg13g2_fill_2 FILLER_0_33_590 ();
 sg13g2_fill_4 FILLER_0_33_597 ();
 sg13g2_fill_8 FILLER_0_33_605 ();
 sg13g2_fill_2 FILLER_0_33_613 ();
 sg13g2_fill_1 FILLER_0_33_615 ();
 sg13g2_fill_2 FILLER_0_33_624 ();
 sg13g2_fill_1 FILLER_0_33_626 ();
 sg13g2_fill_4 FILLER_0_33_632 ();
 sg13g2_fill_2 FILLER_0_33_641 ();
 sg13g2_fill_1 FILLER_0_33_643 ();
 sg13g2_fill_4 FILLER_0_33_648 ();
 sg13g2_fill_8 FILLER_0_33_678 ();
 sg13g2_fill_4 FILLER_0_33_686 ();
 sg13g2_fill_8 FILLER_0_33_695 ();
 sg13g2_fill_1 FILLER_0_33_703 ();
 sg13g2_fill_4 FILLER_0_33_709 ();
 sg13g2_fill_1 FILLER_0_33_713 ();
 sg13g2_fill_4 FILLER_0_33_740 ();
 sg13g2_fill_2 FILLER_0_33_744 ();
 sg13g2_fill_1 FILLER_0_33_746 ();
 sg13g2_fill_4 FILLER_0_33_773 ();
 sg13g2_fill_1 FILLER_0_33_777 ();
 sg13g2_fill_2 FILLER_0_33_783 ();
 sg13g2_fill_4 FILLER_0_33_790 ();
 sg13g2_fill_4 FILLER_0_33_815 ();
 sg13g2_fill_1 FILLER_0_33_819 ();
 sg13g2_fill_2 FILLER_0_33_846 ();
 sg13g2_fill_8 FILLER_0_33_852 ();
 sg13g2_fill_4 FILLER_0_33_860 ();
 sg13g2_fill_2 FILLER_0_33_864 ();
 sg13g2_fill_2 FILLER_0_33_871 ();
 sg13g2_fill_8 FILLER_0_33_877 ();
 sg13g2_fill_8 FILLER_0_33_885 ();
 sg13g2_fill_4 FILLER_0_33_893 ();
 sg13g2_fill_1 FILLER_0_33_897 ();
 sg13g2_fill_4 FILLER_0_33_903 ();
 sg13g2_fill_1 FILLER_0_33_907 ();
 sg13g2_fill_2 FILLER_0_33_912 ();
 sg13g2_fill_8 FILLER_0_33_919 ();
 sg13g2_fill_8 FILLER_0_33_932 ();
 sg13g2_fill_2 FILLER_0_33_944 ();
 sg13g2_fill_4 FILLER_0_33_972 ();
 sg13g2_fill_2 FILLER_0_33_976 ();
 sg13g2_fill_1 FILLER_0_33_978 ();
 sg13g2_fill_2 FILLER_0_33_984 ();
 sg13g2_fill_8 FILLER_0_33_991 ();
 sg13g2_fill_4 FILLER_0_33_999 ();
 sg13g2_fill_2 FILLER_0_33_1003 ();
 sg13g2_fill_2 FILLER_0_33_1010 ();
 sg13g2_fill_8 FILLER_0_33_1016 ();
 sg13g2_fill_8 FILLER_0_33_1024 ();
 sg13g2_fill_2 FILLER_0_33_1032 ();
 sg13g2_fill_1 FILLER_0_33_1034 ();
 sg13g2_fill_2 FILLER_0_33_1056 ();
 sg13g2_fill_8 FILLER_0_33_1079 ();
 sg13g2_fill_8 FILLER_0_33_1087 ();
 sg13g2_fill_4 FILLER_0_33_1095 ();
 sg13g2_fill_8 FILLER_0_33_1103 ();
 sg13g2_fill_8 FILLER_0_33_1111 ();
 sg13g2_fill_8 FILLER_0_33_1119 ();
 sg13g2_fill_1 FILLER_0_33_1127 ();
 sg13g2_fill_2 FILLER_0_33_1132 ();
 sg13g2_fill_2 FILLER_0_33_1140 ();
 sg13g2_fill_8 FILLER_0_33_1146 ();
 sg13g2_fill_1 FILLER_0_33_1154 ();
 sg13g2_fill_2 FILLER_0_33_1162 ();
 sg13g2_fill_2 FILLER_0_33_1169 ();
 sg13g2_fill_1 FILLER_0_33_1171 ();
 sg13g2_fill_2 FILLER_0_33_1180 ();
 sg13g2_fill_2 FILLER_0_33_1187 ();
 sg13g2_fill_4 FILLER_0_33_1196 ();
 sg13g2_fill_2 FILLER_0_33_1207 ();
 sg13g2_fill_2 FILLER_0_33_1214 ();
 sg13g2_fill_1 FILLER_0_33_1216 ();
 sg13g2_fill_4 FILLER_0_33_1223 ();
 sg13g2_fill_8 FILLER_0_33_1231 ();
 sg13g2_fill_8 FILLER_0_33_1239 ();
 sg13g2_fill_8 FILLER_0_33_1247 ();
 sg13g2_fill_8 FILLER_0_33_1255 ();
 sg13g2_fill_4 FILLER_0_33_1263 ();
 sg13g2_fill_2 FILLER_0_33_1267 ();
 sg13g2_fill_2 FILLER_0_33_1295 ();
 sg13g2_fill_8 FILLER_0_34_0 ();
 sg13g2_fill_8 FILLER_0_34_8 ();
 sg13g2_fill_8 FILLER_0_34_16 ();
 sg13g2_fill_8 FILLER_0_34_24 ();
 sg13g2_fill_8 FILLER_0_34_32 ();
 sg13g2_fill_8 FILLER_0_34_40 ();
 sg13g2_fill_8 FILLER_0_34_48 ();
 sg13g2_fill_8 FILLER_0_34_56 ();
 sg13g2_fill_8 FILLER_0_34_64 ();
 sg13g2_fill_8 FILLER_0_34_72 ();
 sg13g2_fill_8 FILLER_0_34_80 ();
 sg13g2_fill_8 FILLER_0_34_88 ();
 sg13g2_fill_8 FILLER_0_34_96 ();
 sg13g2_fill_8 FILLER_0_34_104 ();
 sg13g2_fill_8 FILLER_0_34_112 ();
 sg13g2_fill_8 FILLER_0_34_120 ();
 sg13g2_fill_8 FILLER_0_34_128 ();
 sg13g2_fill_8 FILLER_0_34_136 ();
 sg13g2_fill_8 FILLER_0_34_144 ();
 sg13g2_fill_8 FILLER_0_34_152 ();
 sg13g2_fill_8 FILLER_0_34_160 ();
 sg13g2_fill_8 FILLER_0_34_168 ();
 sg13g2_fill_8 FILLER_0_34_176 ();
 sg13g2_fill_8 FILLER_0_34_184 ();
 sg13g2_fill_8 FILLER_0_34_192 ();
 sg13g2_fill_8 FILLER_0_34_200 ();
 sg13g2_fill_1 FILLER_0_34_208 ();
 sg13g2_fill_2 FILLER_0_34_214 ();
 sg13g2_fill_8 FILLER_0_34_242 ();
 sg13g2_fill_8 FILLER_0_34_250 ();
 sg13g2_fill_4 FILLER_0_34_258 ();
 sg13g2_fill_1 FILLER_0_34_262 ();
 sg13g2_fill_2 FILLER_0_34_268 ();
 sg13g2_fill_1 FILLER_0_34_270 ();
 sg13g2_fill_8 FILLER_0_34_275 ();
 sg13g2_fill_8 FILLER_0_34_283 ();
 sg13g2_fill_8 FILLER_0_34_291 ();
 sg13g2_fill_8 FILLER_0_34_299 ();
 sg13g2_fill_4 FILLER_0_34_307 ();
 sg13g2_fill_4 FILLER_0_34_332 ();
 sg13g2_fill_2 FILLER_0_34_336 ();
 sg13g2_fill_1 FILLER_0_34_338 ();
 sg13g2_fill_2 FILLER_0_34_344 ();
 sg13g2_fill_8 FILLER_0_34_367 ();
 sg13g2_fill_8 FILLER_0_34_375 ();
 sg13g2_fill_8 FILLER_0_34_383 ();
 sg13g2_fill_8 FILLER_0_34_391 ();
 sg13g2_fill_8 FILLER_0_34_399 ();
 sg13g2_fill_4 FILLER_0_34_407 ();
 sg13g2_fill_2 FILLER_0_34_411 ();
 sg13g2_fill_2 FILLER_0_34_418 ();
 sg13g2_fill_2 FILLER_0_34_425 ();
 sg13g2_fill_2 FILLER_0_34_453 ();
 sg13g2_fill_8 FILLER_0_34_476 ();
 sg13g2_fill_8 FILLER_0_34_484 ();
 sg13g2_fill_8 FILLER_0_34_492 ();
 sg13g2_fill_8 FILLER_0_34_500 ();
 sg13g2_fill_2 FILLER_0_34_508 ();
 sg13g2_fill_2 FILLER_0_34_515 ();
 sg13g2_fill_2 FILLER_0_34_521 ();
 sg13g2_fill_1 FILLER_0_34_523 ();
 sg13g2_fill_8 FILLER_0_34_529 ();
 sg13g2_fill_4 FILLER_0_34_537 ();
 sg13g2_fill_2 FILLER_0_34_546 ();
 sg13g2_fill_1 FILLER_0_34_548 ();
 sg13g2_fill_8 FILLER_0_34_553 ();
 sg13g2_fill_4 FILLER_0_34_561 ();
 sg13g2_fill_2 FILLER_0_34_586 ();
 sg13g2_fill_4 FILLER_0_34_595 ();
 sg13g2_fill_2 FILLER_0_34_599 ();
 sg13g2_fill_1 FILLER_0_34_601 ();
 sg13g2_fill_4 FILLER_0_34_609 ();
 sg13g2_fill_2 FILLER_0_34_613 ();
 sg13g2_fill_1 FILLER_0_34_615 ();
 sg13g2_fill_8 FILLER_0_34_628 ();
 sg13g2_fill_2 FILLER_0_34_636 ();
 sg13g2_fill_1 FILLER_0_34_638 ();
 sg13g2_fill_8 FILLER_0_34_665 ();
 sg13g2_fill_8 FILLER_0_34_673 ();
 sg13g2_fill_4 FILLER_0_34_681 ();
 sg13g2_fill_8 FILLER_0_34_690 ();
 sg13g2_fill_4 FILLER_0_34_698 ();
 sg13g2_fill_2 FILLER_0_34_702 ();
 sg13g2_fill_1 FILLER_0_34_704 ();
 sg13g2_fill_2 FILLER_0_34_731 ();
 sg13g2_fill_2 FILLER_0_34_743 ();
 sg13g2_fill_8 FILLER_0_34_749 ();
 sg13g2_fill_4 FILLER_0_34_757 ();
 sg13g2_fill_2 FILLER_0_34_761 ();
 sg13g2_fill_8 FILLER_0_34_768 ();
 sg13g2_fill_8 FILLER_0_34_776 ();
 sg13g2_fill_8 FILLER_0_34_784 ();
 sg13g2_fill_8 FILLER_0_34_792 ();
 sg13g2_fill_1 FILLER_0_34_800 ();
 sg13g2_fill_4 FILLER_0_34_811 ();
 sg13g2_fill_1 FILLER_0_34_815 ();
 sg13g2_fill_8 FILLER_0_34_821 ();
 sg13g2_fill_2 FILLER_0_34_834 ();
 sg13g2_fill_2 FILLER_0_34_840 ();
 sg13g2_fill_1 FILLER_0_34_842 ();
 sg13g2_fill_8 FILLER_0_34_847 ();
 sg13g2_fill_8 FILLER_0_34_855 ();
 sg13g2_fill_8 FILLER_0_34_863 ();
 sg13g2_fill_8 FILLER_0_34_871 ();
 sg13g2_fill_8 FILLER_0_34_879 ();
 sg13g2_fill_4 FILLER_0_34_887 ();
 sg13g2_fill_8 FILLER_0_34_899 ();
 sg13g2_fill_4 FILLER_0_34_907 ();
 sg13g2_fill_2 FILLER_0_34_911 ();
 sg13g2_fill_8 FILLER_0_34_918 ();
 sg13g2_fill_8 FILLER_0_34_926 ();
 sg13g2_fill_8 FILLER_0_34_934 ();
 sg13g2_fill_8 FILLER_0_34_942 ();
 sg13g2_fill_8 FILLER_0_34_950 ();
 sg13g2_fill_8 FILLER_0_34_958 ();
 sg13g2_fill_8 FILLER_0_34_966 ();
 sg13g2_fill_1 FILLER_0_34_974 ();
 sg13g2_fill_8 FILLER_0_34_980 ();
 sg13g2_fill_2 FILLER_0_34_988 ();
 sg13g2_fill_2 FILLER_0_34_995 ();
 sg13g2_fill_8 FILLER_0_34_1001 ();
 sg13g2_fill_8 FILLER_0_34_1009 ();
 sg13g2_fill_8 FILLER_0_34_1017 ();
 sg13g2_fill_8 FILLER_0_34_1025 ();
 sg13g2_fill_8 FILLER_0_34_1033 ();
 sg13g2_fill_8 FILLER_0_34_1041 ();
 sg13g2_fill_8 FILLER_0_34_1049 ();
 sg13g2_fill_4 FILLER_0_34_1057 ();
 sg13g2_fill_2 FILLER_0_34_1061 ();
 sg13g2_fill_8 FILLER_0_34_1067 ();
 sg13g2_fill_2 FILLER_0_34_1075 ();
 sg13g2_fill_8 FILLER_0_34_1082 ();
 sg13g2_fill_4 FILLER_0_34_1090 ();
 sg13g2_fill_2 FILLER_0_34_1099 ();
 sg13g2_fill_4 FILLER_0_34_1105 ();
 sg13g2_fill_8 FILLER_0_34_1115 ();
 sg13g2_fill_8 FILLER_0_34_1123 ();
 sg13g2_fill_2 FILLER_0_34_1131 ();
 sg13g2_fill_2 FILLER_0_34_1138 ();
 sg13g2_fill_2 FILLER_0_34_1145 ();
 sg13g2_fill_1 FILLER_0_34_1147 ();
 sg13g2_fill_2 FILLER_0_34_1156 ();
 sg13g2_fill_1 FILLER_0_34_1158 ();
 sg13g2_fill_2 FILLER_0_34_1165 ();
 sg13g2_fill_1 FILLER_0_34_1167 ();
 sg13g2_fill_2 FILLER_0_34_1173 ();
 sg13g2_fill_1 FILLER_0_34_1175 ();
 sg13g2_fill_2 FILLER_0_34_1180 ();
 sg13g2_fill_1 FILLER_0_34_1182 ();
 sg13g2_fill_8 FILLER_0_34_1191 ();
 sg13g2_fill_8 FILLER_0_34_1199 ();
 sg13g2_fill_8 FILLER_0_34_1207 ();
 sg13g2_fill_2 FILLER_0_34_1215 ();
 sg13g2_fill_2 FILLER_0_34_1222 ();
 sg13g2_fill_8 FILLER_0_34_1230 ();
 sg13g2_fill_8 FILLER_0_34_1238 ();
 sg13g2_fill_8 FILLER_0_34_1246 ();
 sg13g2_fill_2 FILLER_0_34_1254 ();
 sg13g2_fill_2 FILLER_0_34_1260 ();
 sg13g2_fill_4 FILLER_0_34_1272 ();
 sg13g2_fill_2 FILLER_0_34_1276 ();
 sg13g2_fill_1 FILLER_0_34_1278 ();
 sg13g2_fill_8 FILLER_0_34_1287 ();
 sg13g2_fill_2 FILLER_0_34_1295 ();
 sg13g2_fill_8 FILLER_0_35_0 ();
 sg13g2_fill_8 FILLER_0_35_8 ();
 sg13g2_fill_8 FILLER_0_35_16 ();
 sg13g2_fill_8 FILLER_0_35_24 ();
 sg13g2_fill_8 FILLER_0_35_32 ();
 sg13g2_fill_8 FILLER_0_35_40 ();
 sg13g2_fill_8 FILLER_0_35_48 ();
 sg13g2_fill_8 FILLER_0_35_56 ();
 sg13g2_fill_8 FILLER_0_35_64 ();
 sg13g2_fill_8 FILLER_0_35_72 ();
 sg13g2_fill_8 FILLER_0_35_80 ();
 sg13g2_fill_8 FILLER_0_35_88 ();
 sg13g2_fill_8 FILLER_0_35_96 ();
 sg13g2_fill_8 FILLER_0_35_104 ();
 sg13g2_fill_8 FILLER_0_35_112 ();
 sg13g2_fill_8 FILLER_0_35_120 ();
 sg13g2_fill_8 FILLER_0_35_128 ();
 sg13g2_fill_8 FILLER_0_35_136 ();
 sg13g2_fill_8 FILLER_0_35_144 ();
 sg13g2_fill_8 FILLER_0_35_152 ();
 sg13g2_fill_8 FILLER_0_35_160 ();
 sg13g2_fill_8 FILLER_0_35_168 ();
 sg13g2_fill_8 FILLER_0_35_176 ();
 sg13g2_fill_8 FILLER_0_35_184 ();
 sg13g2_fill_8 FILLER_0_35_192 ();
 sg13g2_fill_8 FILLER_0_35_200 ();
 sg13g2_fill_8 FILLER_0_35_208 ();
 sg13g2_fill_2 FILLER_0_35_216 ();
 sg13g2_fill_1 FILLER_0_35_218 ();
 sg13g2_fill_2 FILLER_0_35_245 ();
 sg13g2_fill_2 FILLER_0_35_251 ();
 sg13g2_fill_1 FILLER_0_35_253 ();
 sg13g2_fill_8 FILLER_0_35_259 ();
 sg13g2_fill_8 FILLER_0_35_267 ();
 sg13g2_fill_4 FILLER_0_35_275 ();
 sg13g2_fill_2 FILLER_0_35_279 ();
 sg13g2_fill_1 FILLER_0_35_281 ();
 sg13g2_fill_4 FILLER_0_35_287 ();
 sg13g2_fill_2 FILLER_0_35_317 ();
 sg13g2_fill_4 FILLER_0_35_322 ();
 sg13g2_fill_2 FILLER_0_35_326 ();
 sg13g2_fill_2 FILLER_0_35_354 ();
 sg13g2_fill_1 FILLER_0_35_356 ();
 sg13g2_fill_4 FILLER_0_35_367 ();
 sg13g2_fill_1 FILLER_0_35_371 ();
 sg13g2_fill_8 FILLER_0_35_377 ();
 sg13g2_fill_4 FILLER_0_35_385 ();
 sg13g2_fill_2 FILLER_0_35_389 ();
 sg13g2_fill_1 FILLER_0_35_391 ();
 sg13g2_fill_2 FILLER_0_35_397 ();
 sg13g2_fill_8 FILLER_0_35_403 ();
 sg13g2_fill_8 FILLER_0_35_411 ();
 sg13g2_fill_8 FILLER_0_35_419 ();
 sg13g2_fill_8 FILLER_0_35_427 ();
 sg13g2_fill_8 FILLER_0_35_435 ();
 sg13g2_fill_8 FILLER_0_35_443 ();
 sg13g2_fill_8 FILLER_0_35_451 ();
 sg13g2_fill_8 FILLER_0_35_459 ();
 sg13g2_fill_8 FILLER_0_35_467 ();
 sg13g2_fill_8 FILLER_0_35_475 ();
 sg13g2_fill_8 FILLER_0_35_483 ();
 sg13g2_fill_8 FILLER_0_35_491 ();
 sg13g2_fill_4 FILLER_0_35_499 ();
 sg13g2_fill_2 FILLER_0_35_503 ();
 sg13g2_fill_1 FILLER_0_35_505 ();
 sg13g2_fill_4 FILLER_0_35_532 ();
 sg13g2_fill_2 FILLER_0_35_536 ();
 sg13g2_fill_1 FILLER_0_35_538 ();
 sg13g2_fill_8 FILLER_0_35_565 ();
 sg13g2_fill_8 FILLER_0_35_573 ();
 sg13g2_fill_8 FILLER_0_35_581 ();
 sg13g2_fill_8 FILLER_0_35_589 ();
 sg13g2_fill_2 FILLER_0_35_597 ();
 sg13g2_fill_1 FILLER_0_35_599 ();
 sg13g2_fill_8 FILLER_0_35_608 ();
 sg13g2_fill_8 FILLER_0_35_616 ();
 sg13g2_fill_8 FILLER_0_35_624 ();
 sg13g2_fill_4 FILLER_0_35_632 ();
 sg13g2_fill_2 FILLER_0_35_636 ();
 sg13g2_fill_1 FILLER_0_35_638 ();
 sg13g2_fill_2 FILLER_0_35_644 ();
 sg13g2_fill_4 FILLER_0_35_667 ();
 sg13g2_fill_2 FILLER_0_35_675 ();
 sg13g2_fill_8 FILLER_0_35_682 ();
 sg13g2_fill_4 FILLER_0_35_690 ();
 sg13g2_fill_1 FILLER_0_35_694 ();
 sg13g2_fill_2 FILLER_0_35_700 ();
 sg13g2_fill_8 FILLER_0_35_710 ();
 sg13g2_fill_8 FILLER_0_35_718 ();
 sg13g2_fill_8 FILLER_0_35_726 ();
 sg13g2_fill_8 FILLER_0_35_734 ();
 sg13g2_fill_8 FILLER_0_35_742 ();
 sg13g2_fill_8 FILLER_0_35_750 ();
 sg13g2_fill_2 FILLER_0_35_758 ();
 sg13g2_fill_8 FILLER_0_35_765 ();
 sg13g2_fill_8 FILLER_0_35_773 ();
 sg13g2_fill_8 FILLER_0_35_781 ();
 sg13g2_fill_4 FILLER_0_35_789 ();
 sg13g2_fill_1 FILLER_0_35_793 ();
 sg13g2_fill_8 FILLER_0_35_799 ();
 sg13g2_fill_1 FILLER_0_35_807 ();
 sg13g2_fill_4 FILLER_0_35_813 ();
 sg13g2_fill_1 FILLER_0_35_817 ();
 sg13g2_fill_2 FILLER_0_35_844 ();
 sg13g2_fill_8 FILLER_0_35_851 ();
 sg13g2_fill_8 FILLER_0_35_859 ();
 sg13g2_fill_8 FILLER_0_35_867 ();
 sg13g2_fill_4 FILLER_0_35_875 ();
 sg13g2_fill_2 FILLER_0_35_879 ();
 sg13g2_fill_2 FILLER_0_35_907 ();
 sg13g2_fill_4 FILLER_0_35_930 ();
 sg13g2_fill_8 FILLER_0_35_960 ();
 sg13g2_fill_4 FILLER_0_35_968 ();
 sg13g2_fill_1 FILLER_0_35_972 ();
 sg13g2_fill_8 FILLER_0_35_981 ();
 sg13g2_fill_8 FILLER_0_35_989 ();
 sg13g2_fill_8 FILLER_0_35_997 ();
 sg13g2_fill_8 FILLER_0_35_1005 ();
 sg13g2_fill_8 FILLER_0_35_1013 ();
 sg13g2_fill_8 FILLER_0_35_1021 ();
 sg13g2_fill_4 FILLER_0_35_1029 ();
 sg13g2_fill_2 FILLER_0_35_1033 ();
 sg13g2_fill_1 FILLER_0_35_1035 ();
 sg13g2_fill_8 FILLER_0_35_1041 ();
 sg13g2_fill_1 FILLER_0_35_1049 ();
 sg13g2_fill_2 FILLER_0_35_1053 ();
 sg13g2_fill_8 FILLER_0_35_1060 ();
 sg13g2_fill_8 FILLER_0_35_1068 ();
 sg13g2_fill_2 FILLER_0_35_1076 ();
 sg13g2_fill_8 FILLER_0_35_1086 ();
 sg13g2_fill_8 FILLER_0_35_1094 ();
 sg13g2_fill_8 FILLER_0_35_1102 ();
 sg13g2_fill_8 FILLER_0_35_1110 ();
 sg13g2_fill_4 FILLER_0_35_1118 ();
 sg13g2_fill_2 FILLER_0_35_1122 ();
 sg13g2_fill_4 FILLER_0_35_1129 ();
 sg13g2_fill_1 FILLER_0_35_1133 ();
 sg13g2_fill_2 FILLER_0_35_1140 ();
 sg13g2_fill_8 FILLER_0_35_1147 ();
 sg13g2_fill_4 FILLER_0_35_1155 ();
 sg13g2_fill_8 FILLER_0_35_1167 ();
 sg13g2_fill_1 FILLER_0_35_1175 ();
 sg13g2_fill_2 FILLER_0_35_1184 ();
 sg13g2_fill_8 FILLER_0_35_1194 ();
 sg13g2_fill_8 FILLER_0_35_1202 ();
 sg13g2_fill_8 FILLER_0_35_1210 ();
 sg13g2_fill_2 FILLER_0_35_1218 ();
 sg13g2_fill_1 FILLER_0_35_1220 ();
 sg13g2_fill_2 FILLER_0_35_1224 ();
 sg13g2_fill_8 FILLER_0_35_1232 ();
 sg13g2_fill_8 FILLER_0_35_1240 ();
 sg13g2_fill_8 FILLER_0_35_1248 ();
 sg13g2_fill_4 FILLER_0_35_1256 ();
 sg13g2_fill_2 FILLER_0_35_1265 ();
 sg13g2_fill_8 FILLER_0_35_1272 ();
 sg13g2_fill_8 FILLER_0_35_1280 ();
 sg13g2_fill_8 FILLER_0_35_1288 ();
 sg13g2_fill_1 FILLER_0_35_1296 ();
 sg13g2_fill_8 FILLER_0_36_0 ();
 sg13g2_fill_8 FILLER_0_36_8 ();
 sg13g2_fill_8 FILLER_0_36_16 ();
 sg13g2_fill_8 FILLER_0_36_24 ();
 sg13g2_fill_8 FILLER_0_36_32 ();
 sg13g2_fill_8 FILLER_0_36_40 ();
 sg13g2_fill_8 FILLER_0_36_48 ();
 sg13g2_fill_8 FILLER_0_36_56 ();
 sg13g2_fill_8 FILLER_0_36_64 ();
 sg13g2_fill_8 FILLER_0_36_72 ();
 sg13g2_fill_8 FILLER_0_36_80 ();
 sg13g2_fill_8 FILLER_0_36_88 ();
 sg13g2_fill_8 FILLER_0_36_96 ();
 sg13g2_fill_8 FILLER_0_36_104 ();
 sg13g2_fill_8 FILLER_0_36_112 ();
 sg13g2_fill_8 FILLER_0_36_120 ();
 sg13g2_fill_8 FILLER_0_36_128 ();
 sg13g2_fill_8 FILLER_0_36_136 ();
 sg13g2_fill_8 FILLER_0_36_144 ();
 sg13g2_fill_8 FILLER_0_36_152 ();
 sg13g2_fill_8 FILLER_0_36_160 ();
 sg13g2_fill_8 FILLER_0_36_168 ();
 sg13g2_fill_8 FILLER_0_36_176 ();
 sg13g2_fill_8 FILLER_0_36_184 ();
 sg13g2_fill_8 FILLER_0_36_192 ();
 sg13g2_fill_8 FILLER_0_36_200 ();
 sg13g2_fill_8 FILLER_0_36_208 ();
 sg13g2_fill_8 FILLER_0_36_216 ();
 sg13g2_fill_8 FILLER_0_36_224 ();
 sg13g2_fill_8 FILLER_0_36_232 ();
 sg13g2_fill_8 FILLER_0_36_240 ();
 sg13g2_fill_8 FILLER_0_36_248 ();
 sg13g2_fill_4 FILLER_0_36_256 ();
 sg13g2_fill_2 FILLER_0_36_260 ();
 sg13g2_fill_1 FILLER_0_36_262 ();
 sg13g2_fill_4 FILLER_0_36_268 ();
 sg13g2_fill_8 FILLER_0_36_276 ();
 sg13g2_fill_8 FILLER_0_36_284 ();
 sg13g2_fill_1 FILLER_0_36_292 ();
 sg13g2_fill_8 FILLER_0_36_297 ();
 sg13g2_fill_8 FILLER_0_36_305 ();
 sg13g2_fill_8 FILLER_0_36_313 ();
 sg13g2_fill_8 FILLER_0_36_321 ();
 sg13g2_fill_2 FILLER_0_36_334 ();
 sg13g2_fill_2 FILLER_0_36_340 ();
 sg13g2_fill_8 FILLER_0_36_368 ();
 sg13g2_fill_2 FILLER_0_36_381 ();
 sg13g2_fill_8 FILLER_0_36_409 ();
 sg13g2_fill_8 FILLER_0_36_417 ();
 sg13g2_fill_4 FILLER_0_36_425 ();
 sg13g2_fill_8 FILLER_0_36_437 ();
 sg13g2_fill_8 FILLER_0_36_445 ();
 sg13g2_fill_2 FILLER_0_36_453 ();
 sg13g2_fill_2 FILLER_0_36_463 ();
 sg13g2_fill_8 FILLER_0_36_470 ();
 sg13g2_fill_8 FILLER_0_36_478 ();
 sg13g2_fill_4 FILLER_0_36_486 ();
 sg13g2_fill_2 FILLER_0_36_490 ();
 sg13g2_fill_1 FILLER_0_36_492 ();
 sg13g2_fill_2 FILLER_0_36_498 ();
 sg13g2_fill_1 FILLER_0_36_500 ();
 sg13g2_fill_8 FILLER_0_36_505 ();
 sg13g2_fill_8 FILLER_0_36_513 ();
 sg13g2_fill_8 FILLER_0_36_521 ();
 sg13g2_fill_8 FILLER_0_36_533 ();
 sg13g2_fill_8 FILLER_0_36_541 ();
 sg13g2_fill_2 FILLER_0_36_549 ();
 sg13g2_fill_4 FILLER_0_36_556 ();
 sg13g2_fill_2 FILLER_0_36_560 ();
 sg13g2_fill_1 FILLER_0_36_562 ();
 sg13g2_fill_8 FILLER_0_36_567 ();
 sg13g2_fill_8 FILLER_0_36_575 ();
 sg13g2_fill_4 FILLER_0_36_583 ();
 sg13g2_fill_2 FILLER_0_36_587 ();
 sg13g2_fill_2 FILLER_0_36_594 ();
 sg13g2_fill_1 FILLER_0_36_596 ();
 sg13g2_fill_8 FILLER_0_36_602 ();
 sg13g2_fill_8 FILLER_0_36_610 ();
 sg13g2_fill_8 FILLER_0_36_618 ();
 sg13g2_fill_4 FILLER_0_36_626 ();
 sg13g2_fill_1 FILLER_0_36_630 ();
 sg13g2_fill_2 FILLER_0_36_636 ();
 sg13g2_fill_8 FILLER_0_36_642 ();
 sg13g2_fill_4 FILLER_0_36_650 ();
 sg13g2_fill_2 FILLER_0_36_654 ();
 sg13g2_fill_1 FILLER_0_36_656 ();
 sg13g2_fill_8 FILLER_0_36_678 ();
 sg13g2_fill_8 FILLER_0_36_686 ();
 sg13g2_fill_4 FILLER_0_36_694 ();
 sg13g2_fill_2 FILLER_0_36_698 ();
 sg13g2_fill_4 FILLER_0_36_705 ();
 sg13g2_fill_4 FILLER_0_36_714 ();
 sg13g2_fill_2 FILLER_0_36_722 ();
 sg13g2_fill_2 FILLER_0_36_728 ();
 sg13g2_fill_2 FILLER_0_36_735 ();
 sg13g2_fill_2 FILLER_0_36_741 ();
 sg13g2_fill_4 FILLER_0_36_748 ();
 sg13g2_fill_1 FILLER_0_36_752 ();
 sg13g2_fill_2 FILLER_0_36_761 ();
 sg13g2_fill_2 FILLER_0_36_768 ();
 sg13g2_fill_4 FILLER_0_36_778 ();
 sg13g2_fill_1 FILLER_0_36_782 ();
 sg13g2_fill_2 FILLER_0_36_787 ();
 sg13g2_fill_8 FILLER_0_36_793 ();
 sg13g2_fill_8 FILLER_0_36_801 ();
 sg13g2_fill_4 FILLER_0_36_809 ();
 sg13g2_fill_8 FILLER_0_36_818 ();
 sg13g2_fill_8 FILLER_0_36_826 ();
 sg13g2_fill_4 FILLER_0_36_834 ();
 sg13g2_fill_1 FILLER_0_36_838 ();
 sg13g2_fill_4 FILLER_0_36_844 ();
 sg13g2_fill_2 FILLER_0_36_848 ();
 sg13g2_fill_8 FILLER_0_36_858 ();
 sg13g2_fill_8 FILLER_0_36_866 ();
 sg13g2_fill_2 FILLER_0_36_874 ();
 sg13g2_fill_2 FILLER_0_36_902 ();
 sg13g2_fill_8 FILLER_0_36_925 ();
 sg13g2_fill_2 FILLER_0_36_933 ();
 sg13g2_fill_2 FILLER_0_36_940 ();
 sg13g2_fill_8 FILLER_0_36_946 ();
 sg13g2_fill_8 FILLER_0_36_954 ();
 sg13g2_fill_8 FILLER_0_36_962 ();
 sg13g2_fill_8 FILLER_0_36_970 ();
 sg13g2_fill_8 FILLER_0_36_978 ();
 sg13g2_fill_2 FILLER_0_36_986 ();
 sg13g2_fill_2 FILLER_0_36_992 ();
 sg13g2_fill_2 FILLER_0_36_998 ();
 sg13g2_fill_2 FILLER_0_36_1004 ();
 sg13g2_fill_1 FILLER_0_36_1006 ();
 sg13g2_fill_4 FILLER_0_36_1033 ();
 sg13g2_fill_8 FILLER_0_36_1058 ();
 sg13g2_fill_4 FILLER_0_36_1066 ();
 sg13g2_fill_2 FILLER_0_36_1070 ();
 sg13g2_fill_8 FILLER_0_36_1077 ();
 sg13g2_fill_8 FILLER_0_36_1085 ();
 sg13g2_fill_8 FILLER_0_36_1093 ();
 sg13g2_fill_4 FILLER_0_36_1101 ();
 sg13g2_fill_2 FILLER_0_36_1113 ();
 sg13g2_fill_4 FILLER_0_36_1120 ();
 sg13g2_fill_2 FILLER_0_36_1124 ();
 sg13g2_fill_2 FILLER_0_36_1130 ();
 sg13g2_fill_1 FILLER_0_36_1132 ();
 sg13g2_fill_4 FILLER_0_36_1138 ();
 sg13g2_fill_2 FILLER_0_36_1142 ();
 sg13g2_fill_1 FILLER_0_36_1144 ();
 sg13g2_fill_8 FILLER_0_36_1150 ();
 sg13g2_fill_8 FILLER_0_36_1158 ();
 sg13g2_fill_8 FILLER_0_36_1166 ();
 sg13g2_fill_8 FILLER_0_36_1174 ();
 sg13g2_fill_8 FILLER_0_36_1182 ();
 sg13g2_fill_4 FILLER_0_36_1190 ();
 sg13g2_fill_2 FILLER_0_36_1194 ();
 sg13g2_fill_8 FILLER_0_36_1201 ();
 sg13g2_fill_2 FILLER_0_36_1209 ();
 sg13g2_fill_1 FILLER_0_36_1211 ();
 sg13g2_fill_2 FILLER_0_36_1220 ();
 sg13g2_fill_2 FILLER_0_36_1226 ();
 sg13g2_fill_2 FILLER_0_36_1233 ();
 sg13g2_fill_8 FILLER_0_36_1243 ();
 sg13g2_fill_4 FILLER_0_36_1251 ();
 sg13g2_fill_2 FILLER_0_36_1255 ();
 sg13g2_fill_1 FILLER_0_36_1257 ();
 sg13g2_fill_8 FILLER_0_36_1284 ();
 sg13g2_fill_4 FILLER_0_36_1292 ();
 sg13g2_fill_1 FILLER_0_36_1296 ();
 sg13g2_fill_8 FILLER_0_37_0 ();
 sg13g2_fill_8 FILLER_0_37_8 ();
 sg13g2_fill_8 FILLER_0_37_16 ();
 sg13g2_fill_8 FILLER_0_37_24 ();
 sg13g2_fill_8 FILLER_0_37_32 ();
 sg13g2_fill_8 FILLER_0_37_40 ();
 sg13g2_fill_8 FILLER_0_37_48 ();
 sg13g2_fill_8 FILLER_0_37_56 ();
 sg13g2_fill_8 FILLER_0_37_64 ();
 sg13g2_fill_8 FILLER_0_37_72 ();
 sg13g2_fill_8 FILLER_0_37_80 ();
 sg13g2_fill_8 FILLER_0_37_88 ();
 sg13g2_fill_8 FILLER_0_37_96 ();
 sg13g2_fill_8 FILLER_0_37_104 ();
 sg13g2_fill_8 FILLER_0_37_112 ();
 sg13g2_fill_8 FILLER_0_37_120 ();
 sg13g2_fill_8 FILLER_0_37_128 ();
 sg13g2_fill_8 FILLER_0_37_136 ();
 sg13g2_fill_8 FILLER_0_37_144 ();
 sg13g2_fill_8 FILLER_0_37_152 ();
 sg13g2_fill_8 FILLER_0_37_160 ();
 sg13g2_fill_8 FILLER_0_37_168 ();
 sg13g2_fill_8 FILLER_0_37_176 ();
 sg13g2_fill_8 FILLER_0_37_184 ();
 sg13g2_fill_8 FILLER_0_37_192 ();
 sg13g2_fill_8 FILLER_0_37_200 ();
 sg13g2_fill_8 FILLER_0_37_208 ();
 sg13g2_fill_8 FILLER_0_37_216 ();
 sg13g2_fill_8 FILLER_0_37_224 ();
 sg13g2_fill_8 FILLER_0_37_232 ();
 sg13g2_fill_8 FILLER_0_37_240 ();
 sg13g2_fill_8 FILLER_0_37_248 ();
 sg13g2_fill_4 FILLER_0_37_256 ();
 sg13g2_fill_1 FILLER_0_37_260 ();
 sg13g2_fill_8 FILLER_0_37_287 ();
 sg13g2_fill_8 FILLER_0_37_295 ();
 sg13g2_fill_8 FILLER_0_37_303 ();
 sg13g2_fill_8 FILLER_0_37_311 ();
 sg13g2_fill_8 FILLER_0_37_319 ();
 sg13g2_fill_8 FILLER_0_37_327 ();
 sg13g2_fill_8 FILLER_0_37_335 ();
 sg13g2_fill_4 FILLER_0_37_343 ();
 sg13g2_fill_2 FILLER_0_37_352 ();
 sg13g2_fill_8 FILLER_0_37_358 ();
 sg13g2_fill_8 FILLER_0_37_366 ();
 sg13g2_fill_1 FILLER_0_37_374 ();
 sg13g2_fill_2 FILLER_0_37_379 ();
 sg13g2_fill_8 FILLER_0_37_407 ();
 sg13g2_fill_8 FILLER_0_37_415 ();
 sg13g2_fill_1 FILLER_0_37_423 ();
 sg13g2_fill_8 FILLER_0_37_429 ();
 sg13g2_fill_4 FILLER_0_37_437 ();
 sg13g2_fill_2 FILLER_0_37_445 ();
 sg13g2_fill_2 FILLER_0_37_455 ();
 sg13g2_fill_2 FILLER_0_37_462 ();
 sg13g2_fill_8 FILLER_0_37_468 ();
 sg13g2_fill_8 FILLER_0_37_476 ();
 sg13g2_fill_8 FILLER_0_37_484 ();
 sg13g2_fill_4 FILLER_0_37_492 ();
 sg13g2_fill_1 FILLER_0_37_496 ();
 sg13g2_fill_2 FILLER_0_37_523 ();
 sg13g2_fill_2 FILLER_0_37_528 ();
 sg13g2_fill_8 FILLER_0_37_535 ();
 sg13g2_fill_8 FILLER_0_37_543 ();
 sg13g2_fill_8 FILLER_0_37_551 ();
 sg13g2_fill_2 FILLER_0_37_559 ();
 sg13g2_fill_2 FILLER_0_37_566 ();
 sg13g2_fill_2 FILLER_0_37_594 ();
 sg13g2_fill_1 FILLER_0_37_596 ();
 sg13g2_fill_8 FILLER_0_37_603 ();
 sg13g2_fill_4 FILLER_0_37_611 ();
 sg13g2_fill_2 FILLER_0_37_615 ();
 sg13g2_fill_2 FILLER_0_37_622 ();
 sg13g2_fill_2 FILLER_0_37_628 ();
 sg13g2_fill_4 FILLER_0_37_656 ();
 sg13g2_fill_2 FILLER_0_37_660 ();
 sg13g2_fill_2 FILLER_0_37_667 ();
 sg13g2_fill_2 FILLER_0_37_673 ();
 sg13g2_fill_8 FILLER_0_37_701 ();
 sg13g2_fill_2 FILLER_0_37_709 ();
 sg13g2_fill_2 FILLER_0_37_716 ();
 sg13g2_fill_1 FILLER_0_37_718 ();
 sg13g2_fill_2 FILLER_0_37_723 ();
 sg13g2_fill_4 FILLER_0_37_731 ();
 sg13g2_fill_4 FILLER_0_37_740 ();
 sg13g2_fill_2 FILLER_0_37_744 ();
 sg13g2_fill_4 FILLER_0_37_752 ();
 sg13g2_fill_2 FILLER_0_37_756 ();
 sg13g2_fill_1 FILLER_0_37_758 ();
 sg13g2_fill_2 FILLER_0_37_764 ();
 sg13g2_fill_8 FILLER_0_37_773 ();
 sg13g2_fill_4 FILLER_0_37_781 ();
 sg13g2_fill_2 FILLER_0_37_785 ();
 sg13g2_fill_1 FILLER_0_37_787 ();
 sg13g2_fill_8 FILLER_0_37_793 ();
 sg13g2_fill_2 FILLER_0_37_801 ();
 sg13g2_fill_8 FILLER_0_37_808 ();
 sg13g2_fill_4 FILLER_0_37_816 ();
 sg13g2_fill_1 FILLER_0_37_820 ();
 sg13g2_fill_4 FILLER_0_37_825 ();
 sg13g2_fill_8 FILLER_0_37_834 ();
 sg13g2_fill_8 FILLER_0_37_842 ();
 sg13g2_fill_8 FILLER_0_37_850 ();
 sg13g2_fill_8 FILLER_0_37_858 ();
 sg13g2_fill_4 FILLER_0_37_866 ();
 sg13g2_fill_2 FILLER_0_37_870 ();
 sg13g2_fill_2 FILLER_0_37_876 ();
 sg13g2_fill_4 FILLER_0_37_883 ();
 sg13g2_fill_2 FILLER_0_37_892 ();
 sg13g2_fill_2 FILLER_0_37_898 ();
 sg13g2_fill_8 FILLER_0_37_926 ();
 sg13g2_fill_8 FILLER_0_37_934 ();
 sg13g2_fill_8 FILLER_0_37_942 ();
 sg13g2_fill_8 FILLER_0_37_950 ();
 sg13g2_fill_8 FILLER_0_37_958 ();
 sg13g2_fill_8 FILLER_0_37_966 ();
 sg13g2_fill_8 FILLER_0_37_974 ();
 sg13g2_fill_2 FILLER_0_37_982 ();
 sg13g2_fill_8 FILLER_0_37_989 ();
 sg13g2_fill_2 FILLER_0_37_1002 ();
 sg13g2_fill_2 FILLER_0_37_1030 ();
 sg13g2_fill_2 FILLER_0_37_1053 ();
 sg13g2_fill_2 FILLER_0_37_1060 ();
 sg13g2_fill_4 FILLER_0_37_1066 ();
 sg13g2_fill_1 FILLER_0_37_1070 ();
 sg13g2_fill_8 FILLER_0_37_1075 ();
 sg13g2_fill_8 FILLER_0_37_1091 ();
 sg13g2_fill_2 FILLER_0_37_1099 ();
 sg13g2_fill_8 FILLER_0_37_1109 ();
 sg13g2_fill_4 FILLER_0_37_1117 ();
 sg13g2_fill_2 FILLER_0_37_1125 ();
 sg13g2_fill_4 FILLER_0_37_1135 ();
 sg13g2_fill_2 FILLER_0_37_1139 ();
 sg13g2_fill_1 FILLER_0_37_1141 ();
 sg13g2_fill_8 FILLER_0_37_1150 ();
 sg13g2_fill_8 FILLER_0_37_1158 ();
 sg13g2_fill_8 FILLER_0_37_1166 ();
 sg13g2_fill_8 FILLER_0_37_1174 ();
 sg13g2_fill_4 FILLER_0_37_1182 ();
 sg13g2_fill_2 FILLER_0_37_1191 ();
 sg13g2_fill_2 FILLER_0_37_1198 ();
 sg13g2_fill_2 FILLER_0_37_1205 ();
 sg13g2_fill_1 FILLER_0_37_1207 ();
 sg13g2_fill_2 FILLER_0_37_1213 ();
 sg13g2_fill_2 FILLER_0_37_1219 ();
 sg13g2_fill_2 FILLER_0_37_1226 ();
 sg13g2_fill_4 FILLER_0_37_1236 ();
 sg13g2_fill_8 FILLER_0_37_1244 ();
 sg13g2_fill_4 FILLER_0_37_1252 ();
 sg13g2_fill_2 FILLER_0_37_1256 ();
 sg13g2_fill_2 FILLER_0_37_1263 ();
 sg13g2_fill_8 FILLER_0_37_1269 ();
 sg13g2_fill_8 FILLER_0_37_1277 ();
 sg13g2_fill_8 FILLER_0_37_1285 ();
 sg13g2_fill_4 FILLER_0_37_1293 ();
 sg13g2_fill_8 FILLER_0_38_0 ();
 sg13g2_fill_8 FILLER_0_38_8 ();
 sg13g2_fill_8 FILLER_0_38_16 ();
 sg13g2_fill_8 FILLER_0_38_24 ();
 sg13g2_fill_8 FILLER_0_38_32 ();
 sg13g2_fill_8 FILLER_0_38_40 ();
 sg13g2_fill_8 FILLER_0_38_48 ();
 sg13g2_fill_8 FILLER_0_38_56 ();
 sg13g2_fill_8 FILLER_0_38_64 ();
 sg13g2_fill_8 FILLER_0_38_72 ();
 sg13g2_fill_8 FILLER_0_38_80 ();
 sg13g2_fill_8 FILLER_0_38_88 ();
 sg13g2_fill_8 FILLER_0_38_96 ();
 sg13g2_fill_8 FILLER_0_38_104 ();
 sg13g2_fill_8 FILLER_0_38_112 ();
 sg13g2_fill_8 FILLER_0_38_120 ();
 sg13g2_fill_8 FILLER_0_38_128 ();
 sg13g2_fill_8 FILLER_0_38_136 ();
 sg13g2_fill_8 FILLER_0_38_144 ();
 sg13g2_fill_8 FILLER_0_38_152 ();
 sg13g2_fill_8 FILLER_0_38_160 ();
 sg13g2_fill_8 FILLER_0_38_168 ();
 sg13g2_fill_8 FILLER_0_38_176 ();
 sg13g2_fill_8 FILLER_0_38_184 ();
 sg13g2_fill_8 FILLER_0_38_192 ();
 sg13g2_fill_8 FILLER_0_38_200 ();
 sg13g2_fill_8 FILLER_0_38_208 ();
 sg13g2_fill_8 FILLER_0_38_216 ();
 sg13g2_fill_8 FILLER_0_38_224 ();
 sg13g2_fill_8 FILLER_0_38_232 ();
 sg13g2_fill_8 FILLER_0_38_240 ();
 sg13g2_fill_2 FILLER_0_38_248 ();
 sg13g2_fill_2 FILLER_0_38_255 ();
 sg13g2_fill_2 FILLER_0_38_262 ();
 sg13g2_fill_8 FILLER_0_38_268 ();
 sg13g2_fill_8 FILLER_0_38_276 ();
 sg13g2_fill_8 FILLER_0_38_284 ();
 sg13g2_fill_8 FILLER_0_38_292 ();
 sg13g2_fill_8 FILLER_0_38_300 ();
 sg13g2_fill_4 FILLER_0_38_308 ();
 sg13g2_fill_1 FILLER_0_38_312 ();
 sg13g2_fill_8 FILLER_0_38_318 ();
 sg13g2_fill_8 FILLER_0_38_330 ();
 sg13g2_fill_8 FILLER_0_38_338 ();
 sg13g2_fill_8 FILLER_0_38_346 ();
 sg13g2_fill_8 FILLER_0_38_354 ();
 sg13g2_fill_8 FILLER_0_38_362 ();
 sg13g2_fill_8 FILLER_0_38_370 ();
 sg13g2_fill_8 FILLER_0_38_378 ();
 sg13g2_fill_8 FILLER_0_38_386 ();
 sg13g2_fill_8 FILLER_0_38_399 ();
 sg13g2_fill_8 FILLER_0_38_407 ();
 sg13g2_fill_8 FILLER_0_38_415 ();
 sg13g2_fill_4 FILLER_0_38_449 ();
 sg13g2_fill_2 FILLER_0_38_453 ();
 sg13g2_fill_1 FILLER_0_38_455 ();
 sg13g2_fill_8 FILLER_0_38_482 ();
 sg13g2_fill_8 FILLER_0_38_490 ();
 sg13g2_fill_8 FILLER_0_38_498 ();
 sg13g2_fill_4 FILLER_0_38_506 ();
 sg13g2_fill_4 FILLER_0_38_531 ();
 sg13g2_fill_1 FILLER_0_38_535 ();
 sg13g2_fill_8 FILLER_0_38_540 ();
 sg13g2_fill_8 FILLER_0_38_552 ();
 sg13g2_fill_8 FILLER_0_38_565 ();
 sg13g2_fill_4 FILLER_0_38_573 ();
 sg13g2_fill_1 FILLER_0_38_577 ();
 sg13g2_fill_8 FILLER_0_38_582 ();
 sg13g2_fill_1 FILLER_0_38_590 ();
 sg13g2_fill_8 FILLER_0_38_594 ();
 sg13g2_fill_2 FILLER_0_38_602 ();
 sg13g2_fill_1 FILLER_0_38_604 ();
 sg13g2_fill_2 FILLER_0_38_631 ();
 sg13g2_fill_1 FILLER_0_38_633 ();
 sg13g2_fill_2 FILLER_0_38_655 ();
 sg13g2_fill_8 FILLER_0_38_661 ();
 sg13g2_fill_8 FILLER_0_38_669 ();
 sg13g2_fill_8 FILLER_0_38_677 ();
 sg13g2_fill_8 FILLER_0_38_685 ();
 sg13g2_fill_2 FILLER_0_38_693 ();
 sg13g2_fill_8 FILLER_0_38_698 ();
 sg13g2_fill_1 FILLER_0_38_706 ();
 sg13g2_fill_2 FILLER_0_38_733 ();
 sg13g2_fill_8 FILLER_0_38_761 ();
 sg13g2_fill_8 FILLER_0_38_769 ();
 sg13g2_fill_2 FILLER_0_38_777 ();
 sg13g2_fill_1 FILLER_0_38_779 ();
 sg13g2_fill_2 FILLER_0_38_806 ();
 sg13g2_fill_2 FILLER_0_38_812 ();
 sg13g2_fill_4 FILLER_0_38_819 ();
 sg13g2_fill_2 FILLER_0_38_823 ();
 sg13g2_fill_2 FILLER_0_38_851 ();
 sg13g2_fill_1 FILLER_0_38_853 ();
 sg13g2_fill_8 FILLER_0_38_859 ();
 sg13g2_fill_8 FILLER_0_38_867 ();
 sg13g2_fill_8 FILLER_0_38_875 ();
 sg13g2_fill_8 FILLER_0_38_887 ();
 sg13g2_fill_2 FILLER_0_38_895 ();
 sg13g2_fill_2 FILLER_0_38_902 ();
 sg13g2_fill_2 FILLER_0_38_909 ();
 sg13g2_fill_1 FILLER_0_38_911 ();
 sg13g2_fill_4 FILLER_0_38_917 ();
 sg13g2_fill_1 FILLER_0_38_921 ();
 sg13g2_fill_8 FILLER_0_38_930 ();
 sg13g2_fill_4 FILLER_0_38_938 ();
 sg13g2_fill_2 FILLER_0_38_946 ();
 sg13g2_fill_2 FILLER_0_38_953 ();
 sg13g2_fill_4 FILLER_0_38_981 ();
 sg13g2_fill_2 FILLER_0_38_985 ();
 sg13g2_fill_1 FILLER_0_38_987 ();
 sg13g2_fill_2 FILLER_0_38_992 ();
 sg13g2_fill_2 FILLER_0_38_999 ();
 sg13g2_fill_8 FILLER_0_38_1009 ();
 sg13g2_fill_2 FILLER_0_38_1022 ();
 sg13g2_fill_2 FILLER_0_38_1032 ();
 sg13g2_fill_4 FILLER_0_38_1039 ();
 sg13g2_fill_1 FILLER_0_38_1043 ();
 sg13g2_fill_2 FILLER_0_38_1070 ();
 sg13g2_fill_8 FILLER_0_38_1077 ();
 sg13g2_fill_8 FILLER_0_38_1085 ();
 sg13g2_fill_8 FILLER_0_38_1093 ();
 sg13g2_fill_2 FILLER_0_38_1109 ();
 sg13g2_fill_8 FILLER_0_38_1118 ();
 sg13g2_fill_8 FILLER_0_38_1126 ();
 sg13g2_fill_8 FILLER_0_38_1134 ();
 sg13g2_fill_2 FILLER_0_38_1142 ();
 sg13g2_fill_8 FILLER_0_38_1151 ();
 sg13g2_fill_1 FILLER_0_38_1159 ();
 sg13g2_fill_8 FILLER_0_38_1166 ();
 sg13g2_fill_8 FILLER_0_38_1174 ();
 sg13g2_fill_8 FILLER_0_38_1182 ();
 sg13g2_fill_2 FILLER_0_38_1195 ();
 sg13g2_fill_8 FILLER_0_38_1201 ();
 sg13g2_fill_2 FILLER_0_38_1209 ();
 sg13g2_fill_2 FILLER_0_38_1219 ();
 sg13g2_fill_2 FILLER_0_38_1224 ();
 sg13g2_fill_8 FILLER_0_38_1231 ();
 sg13g2_fill_8 FILLER_0_38_1239 ();
 sg13g2_fill_4 FILLER_0_38_1247 ();
 sg13g2_fill_2 FILLER_0_38_1251 ();
 sg13g2_fill_2 FILLER_0_38_1259 ();
 sg13g2_fill_8 FILLER_0_38_1265 ();
 sg13g2_fill_4 FILLER_0_38_1273 ();
 sg13g2_fill_1 FILLER_0_38_1277 ();
 sg13g2_fill_8 FILLER_0_38_1286 ();
 sg13g2_fill_2 FILLER_0_38_1294 ();
 sg13g2_fill_1 FILLER_0_38_1296 ();
 sg13g2_fill_8 FILLER_0_39_0 ();
 sg13g2_fill_8 FILLER_0_39_8 ();
 sg13g2_fill_8 FILLER_0_39_16 ();
 sg13g2_fill_8 FILLER_0_39_24 ();
 sg13g2_fill_8 FILLER_0_39_32 ();
 sg13g2_fill_8 FILLER_0_39_40 ();
 sg13g2_fill_8 FILLER_0_39_48 ();
 sg13g2_fill_8 FILLER_0_39_56 ();
 sg13g2_fill_8 FILLER_0_39_64 ();
 sg13g2_fill_8 FILLER_0_39_72 ();
 sg13g2_fill_8 FILLER_0_39_80 ();
 sg13g2_fill_8 FILLER_0_39_88 ();
 sg13g2_fill_8 FILLER_0_39_96 ();
 sg13g2_fill_8 FILLER_0_39_104 ();
 sg13g2_fill_8 FILLER_0_39_112 ();
 sg13g2_fill_8 FILLER_0_39_120 ();
 sg13g2_fill_8 FILLER_0_39_128 ();
 sg13g2_fill_8 FILLER_0_39_136 ();
 sg13g2_fill_8 FILLER_0_39_144 ();
 sg13g2_fill_8 FILLER_0_39_152 ();
 sg13g2_fill_8 FILLER_0_39_160 ();
 sg13g2_fill_8 FILLER_0_39_168 ();
 sg13g2_fill_8 FILLER_0_39_176 ();
 sg13g2_fill_8 FILLER_0_39_184 ();
 sg13g2_fill_8 FILLER_0_39_192 ();
 sg13g2_fill_8 FILLER_0_39_200 ();
 sg13g2_fill_8 FILLER_0_39_208 ();
 sg13g2_fill_8 FILLER_0_39_216 ();
 sg13g2_fill_8 FILLER_0_39_229 ();
 sg13g2_fill_4 FILLER_0_39_241 ();
 sg13g2_fill_1 FILLER_0_39_245 ();
 sg13g2_fill_2 FILLER_0_39_272 ();
 sg13g2_fill_8 FILLER_0_39_295 ();
 sg13g2_fill_4 FILLER_0_39_303 ();
 sg13g2_fill_2 FILLER_0_39_307 ();
 sg13g2_fill_8 FILLER_0_39_335 ();
 sg13g2_fill_8 FILLER_0_39_343 ();
 sg13g2_fill_8 FILLER_0_39_351 ();
 sg13g2_fill_8 FILLER_0_39_359 ();
 sg13g2_fill_1 FILLER_0_39_367 ();
 sg13g2_fill_4 FILLER_0_39_373 ();
 sg13g2_fill_1 FILLER_0_39_377 ();
 sg13g2_fill_4 FILLER_0_39_382 ();
 sg13g2_fill_2 FILLER_0_39_386 ();
 sg13g2_fill_1 FILLER_0_39_388 ();
 sg13g2_fill_4 FILLER_0_39_394 ();
 sg13g2_fill_8 FILLER_0_39_419 ();
 sg13g2_fill_4 FILLER_0_39_427 ();
 sg13g2_fill_2 FILLER_0_39_431 ();
 sg13g2_fill_2 FILLER_0_39_459 ();
 sg13g2_fill_2 FILLER_0_39_466 ();
 sg13g2_fill_4 FILLER_0_39_489 ();
 sg13g2_fill_2 FILLER_0_39_519 ();
 sg13g2_fill_4 FILLER_0_39_542 ();
 sg13g2_fill_2 FILLER_0_39_546 ();
 sg13g2_fill_4 FILLER_0_39_552 ();
 sg13g2_fill_2 FILLER_0_39_556 ();
 sg13g2_fill_1 FILLER_0_39_558 ();
 sg13g2_fill_2 FILLER_0_39_585 ();
 sg13g2_fill_8 FILLER_0_39_591 ();
 sg13g2_fill_8 FILLER_0_39_599 ();
 sg13g2_fill_8 FILLER_0_39_607 ();
 sg13g2_fill_2 FILLER_0_39_623 ();
 sg13g2_fill_4 FILLER_0_39_630 ();
 sg13g2_fill_2 FILLER_0_39_634 ();
 sg13g2_fill_2 FILLER_0_39_640 ();
 sg13g2_fill_8 FILLER_0_39_647 ();
 sg13g2_fill_8 FILLER_0_39_655 ();
 sg13g2_fill_8 FILLER_0_39_663 ();
 sg13g2_fill_4 FILLER_0_39_671 ();
 sg13g2_fill_2 FILLER_0_39_675 ();
 sg13g2_fill_1 FILLER_0_39_677 ();
 sg13g2_fill_2 FILLER_0_39_684 ();
 sg13g2_fill_4 FILLER_0_39_690 ();
 sg13g2_fill_1 FILLER_0_39_694 ();
 sg13g2_fill_2 FILLER_0_39_701 ();
 sg13g2_fill_2 FILLER_0_39_708 ();
 sg13g2_fill_8 FILLER_0_39_715 ();
 sg13g2_fill_4 FILLER_0_39_723 ();
 sg13g2_fill_4 FILLER_0_39_732 ();
 sg13g2_fill_2 FILLER_0_39_736 ();
 sg13g2_fill_8 FILLER_0_39_748 ();
 sg13g2_fill_8 FILLER_0_39_756 ();
 sg13g2_fill_8 FILLER_0_39_764 ();
 sg13g2_fill_8 FILLER_0_39_772 ();
 sg13g2_fill_8 FILLER_0_39_780 ();
 sg13g2_fill_8 FILLER_0_39_788 ();
 sg13g2_fill_8 FILLER_0_39_796 ();
 sg13g2_fill_4 FILLER_0_39_804 ();
 sg13g2_fill_1 FILLER_0_39_808 ();
 sg13g2_fill_2 FILLER_0_39_835 ();
 sg13g2_fill_1 FILLER_0_39_837 ();
 sg13g2_fill_2 FILLER_0_39_859 ();
 sg13g2_fill_8 FILLER_0_39_866 ();
 sg13g2_fill_8 FILLER_0_39_874 ();
 sg13g2_fill_8 FILLER_0_39_882 ();
 sg13g2_fill_4 FILLER_0_39_890 ();
 sg13g2_fill_1 FILLER_0_39_894 ();
 sg13g2_fill_8 FILLER_0_39_900 ();
 sg13g2_fill_2 FILLER_0_39_908 ();
 sg13g2_fill_1 FILLER_0_39_910 ();
 sg13g2_fill_2 FILLER_0_39_916 ();
 sg13g2_fill_8 FILLER_0_39_922 ();
 sg13g2_fill_8 FILLER_0_39_930 ();
 sg13g2_fill_8 FILLER_0_39_938 ();
 sg13g2_fill_4 FILLER_0_39_946 ();
 sg13g2_fill_2 FILLER_0_39_954 ();
 sg13g2_fill_2 FILLER_0_39_961 ();
 sg13g2_fill_8 FILLER_0_39_989 ();
 sg13g2_fill_8 FILLER_0_39_997 ();
 sg13g2_fill_8 FILLER_0_39_1005 ();
 sg13g2_fill_2 FILLER_0_39_1013 ();
 sg13g2_fill_2 FILLER_0_39_1019 ();
 sg13g2_fill_8 FILLER_0_39_1047 ();
 sg13g2_fill_8 FILLER_0_39_1055 ();
 sg13g2_fill_8 FILLER_0_39_1063 ();
 sg13g2_fill_8 FILLER_0_39_1071 ();
 sg13g2_fill_8 FILLER_0_39_1079 ();
 sg13g2_fill_2 FILLER_0_39_1087 ();
 sg13g2_fill_1 FILLER_0_39_1089 ();
 sg13g2_fill_2 FILLER_0_39_1095 ();
 sg13g2_fill_1 FILLER_0_39_1097 ();
 sg13g2_fill_8 FILLER_0_39_1103 ();
 sg13g2_fill_8 FILLER_0_39_1111 ();
 sg13g2_fill_8 FILLER_0_39_1119 ();
 sg13g2_fill_1 FILLER_0_39_1127 ();
 sg13g2_fill_8 FILLER_0_39_1132 ();
 sg13g2_fill_1 FILLER_0_39_1140 ();
 sg13g2_fill_2 FILLER_0_39_1149 ();
 sg13g2_fill_8 FILLER_0_39_1161 ();
 sg13g2_fill_8 FILLER_0_39_1169 ();
 sg13g2_fill_8 FILLER_0_39_1177 ();
 sg13g2_fill_8 FILLER_0_39_1185 ();
 sg13g2_fill_8 FILLER_0_39_1193 ();
 sg13g2_fill_8 FILLER_0_39_1201 ();
 sg13g2_fill_4 FILLER_0_39_1209 ();
 sg13g2_fill_2 FILLER_0_39_1213 ();
 sg13g2_fill_1 FILLER_0_39_1215 ();
 sg13g2_fill_8 FILLER_0_39_1221 ();
 sg13g2_fill_4 FILLER_0_39_1229 ();
 sg13g2_fill_2 FILLER_0_39_1233 ();
 sg13g2_fill_1 FILLER_0_39_1235 ();
 sg13g2_fill_8 FILLER_0_39_1246 ();
 sg13g2_fill_2 FILLER_0_39_1254 ();
 sg13g2_fill_1 FILLER_0_39_1256 ();
 sg13g2_fill_4 FILLER_0_39_1267 ();
 sg13g2_fill_2 FILLER_0_39_1279 ();
 sg13g2_fill_8 FILLER_0_39_1285 ();
 sg13g2_fill_4 FILLER_0_39_1293 ();
 sg13g2_fill_8 FILLER_0_40_0 ();
 sg13g2_fill_8 FILLER_0_40_8 ();
 sg13g2_fill_8 FILLER_0_40_16 ();
 sg13g2_fill_8 FILLER_0_40_24 ();
 sg13g2_fill_8 FILLER_0_40_32 ();
 sg13g2_fill_8 FILLER_0_40_40 ();
 sg13g2_fill_8 FILLER_0_40_48 ();
 sg13g2_fill_8 FILLER_0_40_56 ();
 sg13g2_fill_8 FILLER_0_40_64 ();
 sg13g2_fill_8 FILLER_0_40_72 ();
 sg13g2_fill_8 FILLER_0_40_80 ();
 sg13g2_fill_8 FILLER_0_40_88 ();
 sg13g2_fill_8 FILLER_0_40_96 ();
 sg13g2_fill_8 FILLER_0_40_104 ();
 sg13g2_fill_8 FILLER_0_40_112 ();
 sg13g2_fill_8 FILLER_0_40_120 ();
 sg13g2_fill_8 FILLER_0_40_128 ();
 sg13g2_fill_8 FILLER_0_40_136 ();
 sg13g2_fill_8 FILLER_0_40_144 ();
 sg13g2_fill_8 FILLER_0_40_152 ();
 sg13g2_fill_8 FILLER_0_40_160 ();
 sg13g2_fill_8 FILLER_0_40_168 ();
 sg13g2_fill_8 FILLER_0_40_176 ();
 sg13g2_fill_8 FILLER_0_40_184 ();
 sg13g2_fill_8 FILLER_0_40_192 ();
 sg13g2_fill_4 FILLER_0_40_200 ();
 sg13g2_fill_2 FILLER_0_40_204 ();
 sg13g2_fill_1 FILLER_0_40_206 ();
 sg13g2_fill_4 FILLER_0_40_212 ();
 sg13g2_fill_1 FILLER_0_40_216 ();
 sg13g2_fill_8 FILLER_0_40_243 ();
 sg13g2_fill_8 FILLER_0_40_251 ();
 sg13g2_fill_8 FILLER_0_40_259 ();
 sg13g2_fill_4 FILLER_0_40_267 ();
 sg13g2_fill_2 FILLER_0_40_271 ();
 sg13g2_fill_1 FILLER_0_40_273 ();
 sg13g2_fill_4 FILLER_0_40_295 ();
 sg13g2_fill_1 FILLER_0_40_299 ();
 sg13g2_fill_2 FILLER_0_40_326 ();
 sg13g2_fill_8 FILLER_0_40_349 ();
 sg13g2_fill_8 FILLER_0_40_357 ();
 sg13g2_fill_4 FILLER_0_40_391 ();
 sg13g2_fill_1 FILLER_0_40_395 ();
 sg13g2_fill_4 FILLER_0_40_417 ();
 sg13g2_fill_2 FILLER_0_40_421 ();
 sg13g2_fill_4 FILLER_0_40_431 ();
 sg13g2_fill_2 FILLER_0_40_440 ();
 sg13g2_fill_2 FILLER_0_40_446 ();
 sg13g2_fill_2 FILLER_0_40_469 ();
 sg13g2_fill_1 FILLER_0_40_471 ();
 sg13g2_fill_2 FILLER_0_40_480 ();
 sg13g2_fill_4 FILLER_0_40_486 ();
 sg13g2_fill_2 FILLER_0_40_495 ();
 sg13g2_fill_2 FILLER_0_40_501 ();
 sg13g2_fill_8 FILLER_0_40_529 ();
 sg13g2_fill_4 FILLER_0_40_537 ();
 sg13g2_fill_2 FILLER_0_40_541 ();
 sg13g2_fill_1 FILLER_0_40_543 ();
 sg13g2_fill_8 FILLER_0_40_549 ();
 sg13g2_fill_8 FILLER_0_40_565 ();
 sg13g2_fill_2 FILLER_0_40_578 ();
 sg13g2_fill_2 FILLER_0_40_588 ();
 sg13g2_fill_8 FILLER_0_40_598 ();
 sg13g2_fill_8 FILLER_0_40_611 ();
 sg13g2_fill_8 FILLER_0_40_624 ();
 sg13g2_fill_2 FILLER_0_40_637 ();
 sg13g2_fill_8 FILLER_0_40_665 ();
 sg13g2_fill_8 FILLER_0_40_673 ();
 sg13g2_fill_2 FILLER_0_40_681 ();
 sg13g2_fill_2 FILLER_0_40_688 ();
 sg13g2_fill_8 FILLER_0_40_696 ();
 sg13g2_fill_8 FILLER_0_40_704 ();
 sg13g2_fill_8 FILLER_0_40_712 ();
 sg13g2_fill_1 FILLER_0_40_720 ();
 sg13g2_fill_8 FILLER_0_40_726 ();
 sg13g2_fill_8 FILLER_0_40_734 ();
 sg13g2_fill_8 FILLER_0_40_742 ();
 sg13g2_fill_8 FILLER_0_40_750 ();
 sg13g2_fill_8 FILLER_0_40_758 ();
 sg13g2_fill_8 FILLER_0_40_766 ();
 sg13g2_fill_8 FILLER_0_40_774 ();
 sg13g2_fill_8 FILLER_0_40_782 ();
 sg13g2_fill_2 FILLER_0_40_790 ();
 sg13g2_fill_8 FILLER_0_40_797 ();
 sg13g2_fill_4 FILLER_0_40_805 ();
 sg13g2_fill_2 FILLER_0_40_809 ();
 sg13g2_fill_2 FILLER_0_40_818 ();
 sg13g2_fill_2 FILLER_0_40_824 ();
 sg13g2_fill_2 FILLER_0_40_831 ();
 sg13g2_fill_1 FILLER_0_40_833 ();
 sg13g2_fill_2 FILLER_0_40_838 ();
 sg13g2_fill_8 FILLER_0_40_861 ();
 sg13g2_fill_8 FILLER_0_40_869 ();
 sg13g2_fill_8 FILLER_0_40_877 ();
 sg13g2_fill_4 FILLER_0_40_889 ();
 sg13g2_fill_2 FILLER_0_40_893 ();
 sg13g2_fill_2 FILLER_0_40_916 ();
 sg13g2_fill_8 FILLER_0_40_939 ();
 sg13g2_fill_8 FILLER_0_40_947 ();
 sg13g2_fill_2 FILLER_0_40_960 ();
 sg13g2_fill_1 FILLER_0_40_962 ();
 sg13g2_fill_4 FILLER_0_40_968 ();
 sg13g2_fill_2 FILLER_0_40_972 ();
 sg13g2_fill_1 FILLER_0_40_974 ();
 sg13g2_fill_8 FILLER_0_40_985 ();
 sg13g2_fill_8 FILLER_0_40_993 ();
 sg13g2_fill_8 FILLER_0_40_1001 ();
 sg13g2_fill_8 FILLER_0_40_1009 ();
 sg13g2_fill_8 FILLER_0_40_1017 ();
 sg13g2_fill_4 FILLER_0_40_1025 ();
 sg13g2_fill_2 FILLER_0_40_1029 ();
 sg13g2_fill_8 FILLER_0_40_1036 ();
 sg13g2_fill_8 FILLER_0_40_1044 ();
 sg13g2_fill_8 FILLER_0_40_1052 ();
 sg13g2_fill_4 FILLER_0_40_1060 ();
 sg13g2_fill_2 FILLER_0_40_1064 ();
 sg13g2_fill_1 FILLER_0_40_1066 ();
 sg13g2_fill_2 FILLER_0_40_1075 ();
 sg13g2_fill_2 FILLER_0_40_1084 ();
 sg13g2_fill_2 FILLER_0_40_1096 ();
 sg13g2_fill_8 FILLER_0_40_1102 ();
 sg13g2_fill_4 FILLER_0_40_1110 ();
 sg13g2_fill_1 FILLER_0_40_1114 ();
 sg13g2_fill_4 FILLER_0_40_1120 ();
 sg13g2_fill_4 FILLER_0_40_1130 ();
 sg13g2_fill_2 FILLER_0_40_1139 ();
 sg13g2_fill_1 FILLER_0_40_1141 ();
 sg13g2_fill_4 FILLER_0_40_1146 ();
 sg13g2_fill_2 FILLER_0_40_1160 ();
 sg13g2_fill_8 FILLER_0_40_1166 ();
 sg13g2_fill_2 FILLER_0_40_1174 ();
 sg13g2_fill_8 FILLER_0_40_1180 ();
 sg13g2_fill_8 FILLER_0_40_1188 ();
 sg13g2_fill_1 FILLER_0_40_1196 ();
 sg13g2_fill_4 FILLER_0_40_1201 ();
 sg13g2_fill_2 FILLER_0_40_1205 ();
 sg13g2_fill_2 FILLER_0_40_1212 ();
 sg13g2_fill_2 FILLER_0_40_1219 ();
 sg13g2_fill_2 FILLER_0_40_1225 ();
 sg13g2_fill_4 FILLER_0_40_1230 ();
 sg13g2_fill_2 FILLER_0_40_1234 ();
 sg13g2_fill_8 FILLER_0_40_1241 ();
 sg13g2_fill_2 FILLER_0_40_1253 ();
 sg13g2_fill_2 FILLER_0_40_1260 ();
 sg13g2_fill_8 FILLER_0_40_1288 ();
 sg13g2_fill_1 FILLER_0_40_1296 ();
 sg13g2_fill_8 FILLER_0_41_0 ();
 sg13g2_fill_8 FILLER_0_41_8 ();
 sg13g2_fill_8 FILLER_0_41_16 ();
 sg13g2_fill_8 FILLER_0_41_24 ();
 sg13g2_fill_8 FILLER_0_41_32 ();
 sg13g2_fill_8 FILLER_0_41_40 ();
 sg13g2_fill_8 FILLER_0_41_48 ();
 sg13g2_fill_8 FILLER_0_41_56 ();
 sg13g2_fill_8 FILLER_0_41_64 ();
 sg13g2_fill_8 FILLER_0_41_72 ();
 sg13g2_fill_8 FILLER_0_41_80 ();
 sg13g2_fill_8 FILLER_0_41_88 ();
 sg13g2_fill_8 FILLER_0_41_96 ();
 sg13g2_fill_8 FILLER_0_41_104 ();
 sg13g2_fill_8 FILLER_0_41_112 ();
 sg13g2_fill_8 FILLER_0_41_120 ();
 sg13g2_fill_8 FILLER_0_41_128 ();
 sg13g2_fill_8 FILLER_0_41_136 ();
 sg13g2_fill_8 FILLER_0_41_144 ();
 sg13g2_fill_8 FILLER_0_41_152 ();
 sg13g2_fill_8 FILLER_0_41_160 ();
 sg13g2_fill_8 FILLER_0_41_168 ();
 sg13g2_fill_8 FILLER_0_41_176 ();
 sg13g2_fill_8 FILLER_0_41_184 ();
 sg13g2_fill_8 FILLER_0_41_192 ();
 sg13g2_fill_2 FILLER_0_41_226 ();
 sg13g2_fill_8 FILLER_0_41_249 ();
 sg13g2_fill_2 FILLER_0_41_257 ();
 sg13g2_fill_1 FILLER_0_41_259 ();
 sg13g2_fill_2 FILLER_0_41_286 ();
 sg13g2_fill_8 FILLER_0_41_293 ();
 sg13g2_fill_8 FILLER_0_41_305 ();
 sg13g2_fill_8 FILLER_0_41_313 ();
 sg13g2_fill_4 FILLER_0_41_321 ();
 sg13g2_fill_2 FILLER_0_41_325 ();
 sg13g2_fill_1 FILLER_0_41_327 ();
 sg13g2_fill_8 FILLER_0_41_349 ();
 sg13g2_fill_4 FILLER_0_41_357 ();
 sg13g2_fill_8 FILLER_0_41_366 ();
 sg13g2_fill_4 FILLER_0_41_382 ();
 sg13g2_fill_2 FILLER_0_41_386 ();
 sg13g2_fill_8 FILLER_0_41_414 ();
 sg13g2_fill_8 FILLER_0_41_422 ();
 sg13g2_fill_2 FILLER_0_41_435 ();
 sg13g2_fill_2 FILLER_0_41_442 ();
 sg13g2_fill_2 FILLER_0_41_448 ();
 sg13g2_fill_2 FILLER_0_41_458 ();
 sg13g2_fill_8 FILLER_0_41_465 ();
 sg13g2_fill_8 FILLER_0_41_473 ();
 sg13g2_fill_8 FILLER_0_41_481 ();
 sg13g2_fill_8 FILLER_0_41_489 ();
 sg13g2_fill_4 FILLER_0_41_497 ();
 sg13g2_fill_2 FILLER_0_41_506 ();
 sg13g2_fill_8 FILLER_0_41_512 ();
 sg13g2_fill_8 FILLER_0_41_520 ();
 sg13g2_fill_4 FILLER_0_41_528 ();
 sg13g2_fill_8 FILLER_0_41_537 ();
 sg13g2_fill_1 FILLER_0_41_545 ();
 sg13g2_fill_8 FILLER_0_41_553 ();
 sg13g2_fill_8 FILLER_0_41_561 ();
 sg13g2_fill_8 FILLER_0_41_569 ();
 sg13g2_fill_8 FILLER_0_41_577 ();
 sg13g2_fill_4 FILLER_0_41_585 ();
 sg13g2_fill_2 FILLER_0_41_593 ();
 sg13g2_fill_8 FILLER_0_41_621 ();
 sg13g2_fill_8 FILLER_0_41_629 ();
 sg13g2_fill_1 FILLER_0_41_637 ();
 sg13g2_fill_2 FILLER_0_41_643 ();
 sg13g2_fill_4 FILLER_0_41_650 ();
 sg13g2_fill_2 FILLER_0_41_654 ();
 sg13g2_fill_8 FILLER_0_41_660 ();
 sg13g2_fill_2 FILLER_0_41_694 ();
 sg13g2_fill_1 FILLER_0_41_696 ();
 sg13g2_fill_8 FILLER_0_41_702 ();
 sg13g2_fill_8 FILLER_0_41_710 ();
 sg13g2_fill_8 FILLER_0_41_718 ();
 sg13g2_fill_8 FILLER_0_41_726 ();
 sg13g2_fill_8 FILLER_0_41_734 ();
 sg13g2_fill_4 FILLER_0_41_742 ();
 sg13g2_fill_2 FILLER_0_41_746 ();
 sg13g2_fill_2 FILLER_0_41_774 ();
 sg13g2_fill_8 FILLER_0_41_781 ();
 sg13g2_fill_8 FILLER_0_41_789 ();
 sg13g2_fill_8 FILLER_0_41_797 ();
 sg13g2_fill_8 FILLER_0_41_805 ();
 sg13g2_fill_8 FILLER_0_41_813 ();
 sg13g2_fill_4 FILLER_0_41_821 ();
 sg13g2_fill_2 FILLER_0_41_825 ();
 sg13g2_fill_1 FILLER_0_41_827 ();
 sg13g2_fill_2 FILLER_0_41_833 ();
 sg13g2_fill_1 FILLER_0_41_835 ();
 sg13g2_fill_4 FILLER_0_41_840 ();
 sg13g2_fill_4 FILLER_0_41_849 ();
 sg13g2_fill_4 FILLER_0_41_879 ();
 sg13g2_fill_1 FILLER_0_41_883 ();
 sg13g2_fill_4 FILLER_0_41_892 ();
 sg13g2_fill_2 FILLER_0_41_896 ();
 sg13g2_fill_4 FILLER_0_41_903 ();
 sg13g2_fill_1 FILLER_0_41_907 ();
 sg13g2_fill_8 FILLER_0_41_912 ();
 sg13g2_fill_2 FILLER_0_41_920 ();
 sg13g2_fill_1 FILLER_0_41_922 ();
 sg13g2_fill_2 FILLER_0_41_928 ();
 sg13g2_fill_2 FILLER_0_41_935 ();
 sg13g2_fill_2 FILLER_0_41_942 ();
 sg13g2_fill_8 FILLER_0_41_948 ();
 sg13g2_fill_8 FILLER_0_41_956 ();
 sg13g2_fill_8 FILLER_0_41_964 ();
 sg13g2_fill_8 FILLER_0_41_972 ();
 sg13g2_fill_8 FILLER_0_41_980 ();
 sg13g2_fill_8 FILLER_0_41_988 ();
 sg13g2_fill_8 FILLER_0_41_996 ();
 sg13g2_fill_2 FILLER_0_41_1004 ();
 sg13g2_fill_8 FILLER_0_41_1012 ();
 sg13g2_fill_2 FILLER_0_41_1020 ();
 sg13g2_fill_1 FILLER_0_41_1022 ();
 sg13g2_fill_8 FILLER_0_41_1031 ();
 sg13g2_fill_8 FILLER_0_41_1039 ();
 sg13g2_fill_8 FILLER_0_41_1047 ();
 sg13g2_fill_8 FILLER_0_41_1055 ();
 sg13g2_fill_8 FILLER_0_41_1063 ();
 sg13g2_fill_4 FILLER_0_41_1076 ();
 sg13g2_fill_2 FILLER_0_41_1080 ();
 sg13g2_fill_8 FILLER_0_41_1089 ();
 sg13g2_fill_2 FILLER_0_41_1097 ();
 sg13g2_fill_8 FILLER_0_41_1104 ();
 sg13g2_fill_4 FILLER_0_41_1112 ();
 sg13g2_fill_2 FILLER_0_41_1116 ();
 sg13g2_fill_8 FILLER_0_41_1126 ();
 sg13g2_fill_8 FILLER_0_41_1134 ();
 sg13g2_fill_8 FILLER_0_41_1142 ();
 sg13g2_fill_1 FILLER_0_41_1150 ();
 sg13g2_fill_4 FILLER_0_41_1155 ();
 sg13g2_fill_2 FILLER_0_41_1159 ();
 sg13g2_fill_1 FILLER_0_41_1161 ();
 sg13g2_fill_2 FILLER_0_41_1167 ();
 sg13g2_fill_2 FILLER_0_41_1174 ();
 sg13g2_fill_1 FILLER_0_41_1176 ();
 sg13g2_fill_8 FILLER_0_41_1182 ();
 sg13g2_fill_4 FILLER_0_41_1190 ();
 sg13g2_fill_2 FILLER_0_41_1194 ();
 sg13g2_fill_8 FILLER_0_41_1201 ();
 sg13g2_fill_4 FILLER_0_41_1209 ();
 sg13g2_fill_2 FILLER_0_41_1213 ();
 sg13g2_fill_2 FILLER_0_41_1223 ();
 sg13g2_fill_4 FILLER_0_41_1231 ();
 sg13g2_fill_1 FILLER_0_41_1235 ();
 sg13g2_fill_8 FILLER_0_41_1244 ();
 sg13g2_fill_8 FILLER_0_41_1252 ();
 sg13g2_fill_8 FILLER_0_41_1260 ();
 sg13g2_fill_8 FILLER_0_41_1268 ();
 sg13g2_fill_1 FILLER_0_41_1276 ();
 sg13g2_fill_2 FILLER_0_41_1281 ();
 sg13g2_fill_8 FILLER_0_41_1287 ();
 sg13g2_fill_2 FILLER_0_41_1295 ();
 sg13g2_fill_8 FILLER_0_42_0 ();
 sg13g2_fill_8 FILLER_0_42_8 ();
 sg13g2_fill_8 FILLER_0_42_16 ();
 sg13g2_fill_8 FILLER_0_42_24 ();
 sg13g2_fill_8 FILLER_0_42_32 ();
 sg13g2_fill_8 FILLER_0_42_40 ();
 sg13g2_fill_8 FILLER_0_42_48 ();
 sg13g2_fill_8 FILLER_0_42_56 ();
 sg13g2_fill_8 FILLER_0_42_64 ();
 sg13g2_fill_8 FILLER_0_42_72 ();
 sg13g2_fill_8 FILLER_0_42_80 ();
 sg13g2_fill_8 FILLER_0_42_88 ();
 sg13g2_fill_8 FILLER_0_42_96 ();
 sg13g2_fill_8 FILLER_0_42_104 ();
 sg13g2_fill_8 FILLER_0_42_112 ();
 sg13g2_fill_8 FILLER_0_42_120 ();
 sg13g2_fill_8 FILLER_0_42_128 ();
 sg13g2_fill_8 FILLER_0_42_136 ();
 sg13g2_fill_8 FILLER_0_42_144 ();
 sg13g2_fill_8 FILLER_0_42_152 ();
 sg13g2_fill_8 FILLER_0_42_160 ();
 sg13g2_fill_8 FILLER_0_42_168 ();
 sg13g2_fill_8 FILLER_0_42_176 ();
 sg13g2_fill_8 FILLER_0_42_184 ();
 sg13g2_fill_8 FILLER_0_42_192 ();
 sg13g2_fill_8 FILLER_0_42_200 ();
 sg13g2_fill_8 FILLER_0_42_208 ();
 sg13g2_fill_2 FILLER_0_42_216 ();
 sg13g2_fill_4 FILLER_0_42_222 ();
 sg13g2_fill_2 FILLER_0_42_226 ();
 sg13g2_fill_8 FILLER_0_42_249 ();
 sg13g2_fill_1 FILLER_0_42_257 ();
 sg13g2_fill_2 FILLER_0_42_284 ();
 sg13g2_fill_4 FILLER_0_42_290 ();
 sg13g2_fill_1 FILLER_0_42_294 ();
 sg13g2_fill_2 FILLER_0_42_300 ();
 sg13g2_fill_2 FILLER_0_42_328 ();
 sg13g2_fill_2 FILLER_0_42_356 ();
 sg13g2_fill_8 FILLER_0_42_366 ();
 sg13g2_fill_8 FILLER_0_42_379 ();
 sg13g2_fill_4 FILLER_0_42_387 ();
 sg13g2_fill_1 FILLER_0_42_391 ();
 sg13g2_fill_2 FILLER_0_42_397 ();
 sg13g2_fill_2 FILLER_0_42_403 ();
 sg13g2_fill_1 FILLER_0_42_405 ();
 sg13g2_fill_4 FILLER_0_42_411 ();
 sg13g2_fill_2 FILLER_0_42_415 ();
 sg13g2_fill_1 FILLER_0_42_417 ();
 sg13g2_fill_8 FILLER_0_42_424 ();
 sg13g2_fill_8 FILLER_0_42_432 ();
 sg13g2_fill_1 FILLER_0_42_440 ();
 sg13g2_fill_2 FILLER_0_42_467 ();
 sg13g2_fill_1 FILLER_0_42_469 ();
 sg13g2_fill_2 FILLER_0_42_476 ();
 sg13g2_fill_1 FILLER_0_42_478 ();
 sg13g2_fill_8 FILLER_0_42_485 ();
 sg13g2_fill_8 FILLER_0_42_493 ();
 sg13g2_fill_8 FILLER_0_42_501 ();
 sg13g2_fill_8 FILLER_0_42_509 ();
 sg13g2_fill_8 FILLER_0_42_517 ();
 sg13g2_fill_2 FILLER_0_42_525 ();
 sg13g2_fill_2 FILLER_0_42_533 ();
 sg13g2_fill_8 FILLER_0_42_540 ();
 sg13g2_fill_4 FILLER_0_42_548 ();
 sg13g2_fill_4 FILLER_0_42_557 ();
 sg13g2_fill_4 FILLER_0_42_566 ();
 sg13g2_fill_2 FILLER_0_42_574 ();
 sg13g2_fill_4 FILLER_0_42_597 ();
 sg13g2_fill_2 FILLER_0_42_601 ();
 sg13g2_fill_2 FILLER_0_42_608 ();
 sg13g2_fill_2 FILLER_0_42_620 ();
 sg13g2_fill_8 FILLER_0_42_627 ();
 sg13g2_fill_8 FILLER_0_42_635 ();
 sg13g2_fill_8 FILLER_0_42_643 ();
 sg13g2_fill_4 FILLER_0_42_651 ();
 sg13g2_fill_2 FILLER_0_42_655 ();
 sg13g2_fill_2 FILLER_0_42_662 ();
 sg13g2_fill_8 FILLER_0_42_670 ();
 sg13g2_fill_1 FILLER_0_42_678 ();
 sg13g2_fill_8 FILLER_0_42_683 ();
 sg13g2_fill_8 FILLER_0_42_691 ();
 sg13g2_fill_1 FILLER_0_42_699 ();
 sg13g2_fill_4 FILLER_0_42_704 ();
 sg13g2_fill_2 FILLER_0_42_708 ();
 sg13g2_fill_4 FILLER_0_42_736 ();
 sg13g2_fill_1 FILLER_0_42_740 ();
 sg13g2_fill_4 FILLER_0_42_746 ();
 sg13g2_fill_2 FILLER_0_42_754 ();
 sg13g2_fill_4 FILLER_0_42_777 ();
 sg13g2_fill_8 FILLER_0_42_785 ();
 sg13g2_fill_8 FILLER_0_42_793 ();
 sg13g2_fill_8 FILLER_0_42_801 ();
 sg13g2_fill_8 FILLER_0_42_809 ();
 sg13g2_fill_4 FILLER_0_42_817 ();
 sg13g2_fill_2 FILLER_0_42_821 ();
 sg13g2_fill_8 FILLER_0_42_849 ();
 sg13g2_fill_4 FILLER_0_42_857 ();
 sg13g2_fill_2 FILLER_0_42_861 ();
 sg13g2_fill_1 FILLER_0_42_863 ();
 sg13g2_fill_4 FILLER_0_42_869 ();
 sg13g2_fill_2 FILLER_0_42_873 ();
 sg13g2_fill_8 FILLER_0_42_879 ();
 sg13g2_fill_1 FILLER_0_42_887 ();
 sg13g2_fill_2 FILLER_0_42_896 ();
 sg13g2_fill_8 FILLER_0_42_924 ();
 sg13g2_fill_1 FILLER_0_42_932 ();
 sg13g2_fill_8 FILLER_0_42_959 ();
 sg13g2_fill_8 FILLER_0_42_967 ();
 sg13g2_fill_8 FILLER_0_42_975 ();
 sg13g2_fill_2 FILLER_0_42_983 ();
 sg13g2_fill_2 FILLER_0_42_988 ();
 sg13g2_fill_4 FILLER_0_42_994 ();
 sg13g2_fill_1 FILLER_0_42_998 ();
 sg13g2_fill_8 FILLER_0_42_1005 ();
 sg13g2_fill_8 FILLER_0_42_1013 ();
 sg13g2_fill_2 FILLER_0_42_1021 ();
 sg13g2_fill_1 FILLER_0_42_1023 ();
 sg13g2_fill_2 FILLER_0_42_1029 ();
 sg13g2_fill_2 FILLER_0_42_1036 ();
 sg13g2_fill_1 FILLER_0_42_1038 ();
 sg13g2_fill_8 FILLER_0_42_1045 ();
 sg13g2_fill_8 FILLER_0_42_1053 ();
 sg13g2_fill_8 FILLER_0_42_1061 ();
 sg13g2_fill_4 FILLER_0_42_1069 ();
 sg13g2_fill_2 FILLER_0_42_1079 ();
 sg13g2_fill_4 FILLER_0_42_1086 ();
 sg13g2_fill_2 FILLER_0_42_1090 ();
 sg13g2_fill_8 FILLER_0_42_1100 ();
 sg13g2_fill_8 FILLER_0_42_1108 ();
 sg13g2_fill_4 FILLER_0_42_1116 ();
 sg13g2_fill_1 FILLER_0_42_1120 ();
 sg13g2_fill_8 FILLER_0_42_1126 ();
 sg13g2_fill_2 FILLER_0_42_1134 ();
 sg13g2_fill_2 FILLER_0_42_1140 ();
 sg13g2_fill_1 FILLER_0_42_1142 ();
 sg13g2_fill_2 FILLER_0_42_1148 ();
 sg13g2_fill_8 FILLER_0_42_1154 ();
 sg13g2_fill_8 FILLER_0_42_1162 ();
 sg13g2_fill_8 FILLER_0_42_1170 ();
 sg13g2_fill_8 FILLER_0_42_1178 ();
 sg13g2_fill_8 FILLER_0_42_1194 ();
 sg13g2_fill_8 FILLER_0_42_1202 ();
 sg13g2_fill_4 FILLER_0_42_1210 ();
 sg13g2_fill_1 FILLER_0_42_1214 ();
 sg13g2_fill_4 FILLER_0_42_1219 ();
 sg13g2_fill_2 FILLER_0_42_1223 ();
 sg13g2_fill_2 FILLER_0_42_1230 ();
 sg13g2_fill_8 FILLER_0_42_1237 ();
 sg13g2_fill_8 FILLER_0_42_1245 ();
 sg13g2_fill_8 FILLER_0_42_1253 ();
 sg13g2_fill_8 FILLER_0_42_1261 ();
 sg13g2_fill_8 FILLER_0_42_1269 ();
 sg13g2_fill_2 FILLER_0_42_1277 ();
 sg13g2_fill_1 FILLER_0_42_1279 ();
 sg13g2_fill_8 FILLER_0_42_1284 ();
 sg13g2_fill_4 FILLER_0_42_1292 ();
 sg13g2_fill_1 FILLER_0_42_1296 ();
 sg13g2_fill_8 FILLER_0_43_0 ();
 sg13g2_fill_8 FILLER_0_43_8 ();
 sg13g2_fill_8 FILLER_0_43_16 ();
 sg13g2_fill_8 FILLER_0_43_24 ();
 sg13g2_fill_8 FILLER_0_43_32 ();
 sg13g2_fill_8 FILLER_0_43_40 ();
 sg13g2_fill_8 FILLER_0_43_48 ();
 sg13g2_fill_8 FILLER_0_43_56 ();
 sg13g2_fill_8 FILLER_0_43_64 ();
 sg13g2_fill_8 FILLER_0_43_72 ();
 sg13g2_fill_8 FILLER_0_43_80 ();
 sg13g2_fill_8 FILLER_0_43_88 ();
 sg13g2_fill_8 FILLER_0_43_96 ();
 sg13g2_fill_8 FILLER_0_43_104 ();
 sg13g2_fill_8 FILLER_0_43_112 ();
 sg13g2_fill_8 FILLER_0_43_120 ();
 sg13g2_fill_8 FILLER_0_43_128 ();
 sg13g2_fill_8 FILLER_0_43_136 ();
 sg13g2_fill_8 FILLER_0_43_144 ();
 sg13g2_fill_8 FILLER_0_43_152 ();
 sg13g2_fill_8 FILLER_0_43_160 ();
 sg13g2_fill_8 FILLER_0_43_168 ();
 sg13g2_fill_8 FILLER_0_43_176 ();
 sg13g2_fill_8 FILLER_0_43_184 ();
 sg13g2_fill_8 FILLER_0_43_192 ();
 sg13g2_fill_8 FILLER_0_43_200 ();
 sg13g2_fill_4 FILLER_0_43_208 ();
 sg13g2_fill_2 FILLER_0_43_212 ();
 sg13g2_fill_2 FILLER_0_43_219 ();
 sg13g2_fill_8 FILLER_0_43_225 ();
 sg13g2_fill_8 FILLER_0_43_233 ();
 sg13g2_fill_8 FILLER_0_43_241 ();
 sg13g2_fill_8 FILLER_0_43_249 ();
 sg13g2_fill_8 FILLER_0_43_257 ();
 sg13g2_fill_4 FILLER_0_43_265 ();
 sg13g2_fill_2 FILLER_0_43_274 ();
 sg13g2_fill_8 FILLER_0_43_280 ();
 sg13g2_fill_4 FILLER_0_43_288 ();
 sg13g2_fill_1 FILLER_0_43_292 ();
 sg13g2_fill_2 FILLER_0_43_298 ();
 sg13g2_fill_8 FILLER_0_43_305 ();
 sg13g2_fill_2 FILLER_0_43_313 ();
 sg13g2_fill_8 FILLER_0_43_319 ();
 sg13g2_fill_4 FILLER_0_43_327 ();
 sg13g2_fill_2 FILLER_0_43_331 ();
 sg13g2_fill_2 FILLER_0_43_338 ();
 sg13g2_fill_1 FILLER_0_43_340 ();
 sg13g2_fill_8 FILLER_0_43_345 ();
 sg13g2_fill_8 FILLER_0_43_353 ();
 sg13g2_fill_8 FILLER_0_43_361 ();
 sg13g2_fill_4 FILLER_0_43_369 ();
 sg13g2_fill_2 FILLER_0_43_373 ();
 sg13g2_fill_1 FILLER_0_43_375 ();
 sg13g2_fill_8 FILLER_0_43_381 ();
 sg13g2_fill_2 FILLER_0_43_389 ();
 sg13g2_fill_8 FILLER_0_43_396 ();
 sg13g2_fill_8 FILLER_0_43_404 ();
 sg13g2_fill_8 FILLER_0_43_412 ();
 sg13g2_fill_8 FILLER_0_43_420 ();
 sg13g2_fill_8 FILLER_0_43_428 ();
 sg13g2_fill_8 FILLER_0_43_436 ();
 sg13g2_fill_8 FILLER_0_43_444 ();
 sg13g2_fill_8 FILLER_0_43_452 ();
 sg13g2_fill_8 FILLER_0_43_460 ();
 sg13g2_fill_4 FILLER_0_43_468 ();
 sg13g2_fill_1 FILLER_0_43_472 ();
 sg13g2_fill_2 FILLER_0_43_485 ();
 sg13g2_fill_8 FILLER_0_43_492 ();
 sg13g2_fill_4 FILLER_0_43_500 ();
 sg13g2_fill_2 FILLER_0_43_504 ();
 sg13g2_fill_1 FILLER_0_43_506 ();
 sg13g2_fill_2 FILLER_0_43_511 ();
 sg13g2_fill_8 FILLER_0_43_518 ();
 sg13g2_fill_8 FILLER_0_43_526 ();
 sg13g2_fill_8 FILLER_0_43_534 ();
 sg13g2_fill_8 FILLER_0_43_542 ();
 sg13g2_fill_8 FILLER_0_43_550 ();
 sg13g2_fill_2 FILLER_0_43_584 ();
 sg13g2_fill_2 FILLER_0_43_589 ();
 sg13g2_fill_8 FILLER_0_43_617 ();
 sg13g2_fill_8 FILLER_0_43_625 ();
 sg13g2_fill_8 FILLER_0_43_633 ();
 sg13g2_fill_8 FILLER_0_43_641 ();
 sg13g2_fill_1 FILLER_0_43_649 ();
 sg13g2_fill_2 FILLER_0_43_655 ();
 sg13g2_fill_8 FILLER_0_43_661 ();
 sg13g2_fill_8 FILLER_0_43_669 ();
 sg13g2_fill_8 FILLER_0_43_677 ();
 sg13g2_fill_8 FILLER_0_43_685 ();
 sg13g2_fill_8 FILLER_0_43_693 ();
 sg13g2_fill_2 FILLER_0_43_706 ();
 sg13g2_fill_4 FILLER_0_43_734 ();
 sg13g2_fill_2 FILLER_0_43_738 ();
 sg13g2_fill_8 FILLER_0_43_766 ();
 sg13g2_fill_2 FILLER_0_43_774 ();
 sg13g2_fill_8 FILLER_0_43_781 ();
 sg13g2_fill_4 FILLER_0_43_789 ();
 sg13g2_fill_1 FILLER_0_43_793 ();
 sg13g2_fill_2 FILLER_0_43_799 ();
 sg13g2_fill_1 FILLER_0_43_801 ();
 sg13g2_fill_8 FILLER_0_43_807 ();
 sg13g2_fill_1 FILLER_0_43_815 ();
 sg13g2_fill_8 FILLER_0_43_820 ();
 sg13g2_fill_8 FILLER_0_43_828 ();
 sg13g2_fill_4 FILLER_0_43_836 ();
 sg13g2_fill_1 FILLER_0_43_840 ();
 sg13g2_fill_8 FILLER_0_43_846 ();
 sg13g2_fill_8 FILLER_0_43_854 ();
 sg13g2_fill_4 FILLER_0_43_862 ();
 sg13g2_fill_1 FILLER_0_43_866 ();
 sg13g2_fill_8 FILLER_0_43_873 ();
 sg13g2_fill_4 FILLER_0_43_881 ();
 sg13g2_fill_1 FILLER_0_43_885 ();
 sg13g2_fill_2 FILLER_0_43_891 ();
 sg13g2_fill_4 FILLER_0_43_897 ();
 sg13g2_fill_2 FILLER_0_43_901 ();
 sg13g2_fill_1 FILLER_0_43_903 ();
 sg13g2_fill_8 FILLER_0_43_911 ();
 sg13g2_fill_2 FILLER_0_43_919 ();
 sg13g2_fill_4 FILLER_0_43_926 ();
 sg13g2_fill_1 FILLER_0_43_930 ();
 sg13g2_fill_2 FILLER_0_43_936 ();
 sg13g2_fill_1 FILLER_0_43_938 ();
 sg13g2_fill_8 FILLER_0_43_944 ();
 sg13g2_fill_8 FILLER_0_43_952 ();
 sg13g2_fill_8 FILLER_0_43_960 ();
 sg13g2_fill_8 FILLER_0_43_968 ();
 sg13g2_fill_2 FILLER_0_43_980 ();
 sg13g2_fill_2 FILLER_0_43_987 ();
 sg13g2_fill_2 FILLER_0_43_993 ();
 sg13g2_fill_1 FILLER_0_43_995 ();
 sg13g2_fill_4 FILLER_0_43_1001 ();
 sg13g2_fill_2 FILLER_0_43_1005 ();
 sg13g2_fill_1 FILLER_0_43_1007 ();
 sg13g2_fill_8 FILLER_0_43_1013 ();
 sg13g2_fill_4 FILLER_0_43_1021 ();
 sg13g2_fill_4 FILLER_0_43_1031 ();
 sg13g2_fill_2 FILLER_0_43_1040 ();
 sg13g2_fill_1 FILLER_0_43_1042 ();
 sg13g2_fill_8 FILLER_0_43_1048 ();
 sg13g2_fill_8 FILLER_0_43_1056 ();
 sg13g2_fill_4 FILLER_0_43_1064 ();
 sg13g2_fill_2 FILLER_0_43_1068 ();
 sg13g2_fill_2 FILLER_0_43_1078 ();
 sg13g2_fill_8 FILLER_0_43_1084 ();
 sg13g2_fill_8 FILLER_0_43_1092 ();
 sg13g2_fill_8 FILLER_0_43_1100 ();
 sg13g2_fill_8 FILLER_0_43_1113 ();
 sg13g2_fill_1 FILLER_0_43_1121 ();
 sg13g2_fill_4 FILLER_0_43_1130 ();
 sg13g2_fill_8 FILLER_0_43_1142 ();
 sg13g2_fill_2 FILLER_0_43_1150 ();
 sg13g2_fill_2 FILLER_0_43_1156 ();
 sg13g2_fill_1 FILLER_0_43_1158 ();
 sg13g2_fill_8 FILLER_0_43_1164 ();
 sg13g2_fill_4 FILLER_0_43_1172 ();
 sg13g2_fill_2 FILLER_0_43_1176 ();
 sg13g2_fill_4 FILLER_0_43_1183 ();
 sg13g2_fill_4 FILLER_0_43_1191 ();
 sg13g2_fill_2 FILLER_0_43_1200 ();
 sg13g2_fill_1 FILLER_0_43_1202 ();
 sg13g2_fill_8 FILLER_0_43_1209 ();
 sg13g2_fill_8 FILLER_0_43_1217 ();
 sg13g2_fill_8 FILLER_0_43_1225 ();
 sg13g2_fill_4 FILLER_0_43_1233 ();
 sg13g2_fill_1 FILLER_0_43_1237 ();
 sg13g2_fill_2 FILLER_0_43_1241 ();
 sg13g2_fill_8 FILLER_0_43_1247 ();
 sg13g2_fill_8 FILLER_0_43_1255 ();
 sg13g2_fill_4 FILLER_0_43_1263 ();
 sg13g2_fill_1 FILLER_0_43_1267 ();
 sg13g2_fill_2 FILLER_0_43_1273 ();
 sg13g2_fill_2 FILLER_0_43_1279 ();
 sg13g2_fill_2 FILLER_0_43_1286 ();
 sg13g2_fill_4 FILLER_0_43_1292 ();
 sg13g2_fill_1 FILLER_0_43_1296 ();
 sg13g2_fill_8 FILLER_0_44_0 ();
 sg13g2_fill_8 FILLER_0_44_8 ();
 sg13g2_fill_8 FILLER_0_44_16 ();
 sg13g2_fill_8 FILLER_0_44_24 ();
 sg13g2_fill_8 FILLER_0_44_32 ();
 sg13g2_fill_8 FILLER_0_44_40 ();
 sg13g2_fill_8 FILLER_0_44_48 ();
 sg13g2_fill_8 FILLER_0_44_56 ();
 sg13g2_fill_8 FILLER_0_44_64 ();
 sg13g2_fill_8 FILLER_0_44_72 ();
 sg13g2_fill_8 FILLER_0_44_80 ();
 sg13g2_fill_8 FILLER_0_44_88 ();
 sg13g2_fill_8 FILLER_0_44_96 ();
 sg13g2_fill_8 FILLER_0_44_104 ();
 sg13g2_fill_8 FILLER_0_44_112 ();
 sg13g2_fill_8 FILLER_0_44_120 ();
 sg13g2_fill_8 FILLER_0_44_128 ();
 sg13g2_fill_8 FILLER_0_44_136 ();
 sg13g2_fill_8 FILLER_0_44_144 ();
 sg13g2_fill_8 FILLER_0_44_152 ();
 sg13g2_fill_8 FILLER_0_44_160 ();
 sg13g2_fill_8 FILLER_0_44_168 ();
 sg13g2_fill_8 FILLER_0_44_176 ();
 sg13g2_fill_8 FILLER_0_44_184 ();
 sg13g2_fill_8 FILLER_0_44_192 ();
 sg13g2_fill_8 FILLER_0_44_200 ();
 sg13g2_fill_2 FILLER_0_44_208 ();
 sg13g2_fill_8 FILLER_0_44_236 ();
 sg13g2_fill_8 FILLER_0_44_244 ();
 sg13g2_fill_8 FILLER_0_44_252 ();
 sg13g2_fill_8 FILLER_0_44_260 ();
 sg13g2_fill_8 FILLER_0_44_268 ();
 sg13g2_fill_8 FILLER_0_44_276 ();
 sg13g2_fill_8 FILLER_0_44_284 ();
 sg13g2_fill_8 FILLER_0_44_292 ();
 sg13g2_fill_8 FILLER_0_44_300 ();
 sg13g2_fill_8 FILLER_0_44_308 ();
 sg13g2_fill_8 FILLER_0_44_316 ();
 sg13g2_fill_8 FILLER_0_44_324 ();
 sg13g2_fill_8 FILLER_0_44_332 ();
 sg13g2_fill_8 FILLER_0_44_340 ();
 sg13g2_fill_8 FILLER_0_44_348 ();
 sg13g2_fill_8 FILLER_0_44_356 ();
 sg13g2_fill_8 FILLER_0_44_364 ();
 sg13g2_fill_8 FILLER_0_44_372 ();
 sg13g2_fill_8 FILLER_0_44_380 ();
 sg13g2_fill_8 FILLER_0_44_388 ();
 sg13g2_fill_8 FILLER_0_44_396 ();
 sg13g2_fill_4 FILLER_0_44_404 ();
 sg13g2_fill_2 FILLER_0_44_408 ();
 sg13g2_fill_8 FILLER_0_44_414 ();
 sg13g2_fill_8 FILLER_0_44_422 ();
 sg13g2_fill_8 FILLER_0_44_430 ();
 sg13g2_fill_8 FILLER_0_44_438 ();
 sg13g2_fill_8 FILLER_0_44_446 ();
 sg13g2_fill_4 FILLER_0_44_454 ();
 sg13g2_fill_2 FILLER_0_44_458 ();
 sg13g2_fill_8 FILLER_0_44_464 ();
 sg13g2_fill_8 FILLER_0_44_472 ();
 sg13g2_fill_4 FILLER_0_44_480 ();
 sg13g2_fill_2 FILLER_0_44_484 ();
 sg13g2_fill_2 FILLER_0_44_512 ();
 sg13g2_fill_1 FILLER_0_44_514 ();
 sg13g2_fill_8 FILLER_0_44_520 ();
 sg13g2_fill_8 FILLER_0_44_528 ();
 sg13g2_fill_4 FILLER_0_44_536 ();
 sg13g2_fill_2 FILLER_0_44_546 ();
 sg13g2_fill_2 FILLER_0_44_552 ();
 sg13g2_fill_2 FILLER_0_44_562 ();
 sg13g2_fill_8 FILLER_0_44_572 ();
 sg13g2_fill_8 FILLER_0_44_580 ();
 sg13g2_fill_1 FILLER_0_44_588 ();
 sg13g2_fill_2 FILLER_0_44_594 ();
 sg13g2_fill_8 FILLER_0_44_600 ();
 sg13g2_fill_2 FILLER_0_44_608 ();
 sg13g2_fill_8 FILLER_0_44_615 ();
 sg13g2_fill_2 FILLER_0_44_623 ();
 sg13g2_fill_1 FILLER_0_44_625 ();
 sg13g2_fill_8 FILLER_0_44_631 ();
 sg13g2_fill_2 FILLER_0_44_639 ();
 sg13g2_fill_2 FILLER_0_44_667 ();
 sg13g2_fill_8 FILLER_0_44_674 ();
 sg13g2_fill_8 FILLER_0_44_682 ();
 sg13g2_fill_8 FILLER_0_44_690 ();
 sg13g2_fill_8 FILLER_0_44_698 ();
 sg13g2_fill_4 FILLER_0_44_706 ();
 sg13g2_fill_1 FILLER_0_44_710 ();
 sg13g2_fill_2 FILLER_0_44_716 ();
 sg13g2_fill_1 FILLER_0_44_718 ();
 sg13g2_fill_8 FILLER_0_44_723 ();
 sg13g2_fill_8 FILLER_0_44_731 ();
 sg13g2_fill_8 FILLER_0_44_739 ();
 sg13g2_fill_8 FILLER_0_44_747 ();
 sg13g2_fill_8 FILLER_0_44_765 ();
 sg13g2_fill_8 FILLER_0_44_773 ();
 sg13g2_fill_8 FILLER_0_44_781 ();
 sg13g2_fill_8 FILLER_0_44_789 ();
 sg13g2_fill_4 FILLER_0_44_797 ();
 sg13g2_fill_1 FILLER_0_44_801 ();
 sg13g2_fill_8 FILLER_0_44_806 ();
 sg13g2_fill_2 FILLER_0_44_814 ();
 sg13g2_fill_1 FILLER_0_44_816 ();
 sg13g2_fill_2 FILLER_0_44_822 ();
 sg13g2_fill_1 FILLER_0_44_824 ();
 sg13g2_fill_2 FILLER_0_44_830 ();
 sg13g2_fill_2 FILLER_0_44_837 ();
 sg13g2_fill_1 FILLER_0_44_839 ();
 sg13g2_fill_8 FILLER_0_44_844 ();
 sg13g2_fill_8 FILLER_0_44_852 ();
 sg13g2_fill_8 FILLER_0_44_860 ();
 sg13g2_fill_8 FILLER_0_44_868 ();
 sg13g2_fill_4 FILLER_0_44_902 ();
 sg13g2_fill_8 FILLER_0_44_911 ();
 sg13g2_fill_8 FILLER_0_44_919 ();
 sg13g2_fill_8 FILLER_0_44_927 ();
 sg13g2_fill_8 FILLER_0_44_935 ();
 sg13g2_fill_8 FILLER_0_44_943 ();
 sg13g2_fill_8 FILLER_0_44_951 ();
 sg13g2_fill_8 FILLER_0_44_959 ();
 sg13g2_fill_8 FILLER_0_44_967 ();
 sg13g2_fill_4 FILLER_0_44_975 ();
 sg13g2_fill_2 FILLER_0_44_979 ();
 sg13g2_fill_1 FILLER_0_44_981 ();
 sg13g2_fill_2 FILLER_0_44_985 ();
 sg13g2_fill_2 FILLER_0_44_992 ();
 sg13g2_fill_2 FILLER_0_44_999 ();
 sg13g2_fill_8 FILLER_0_44_1006 ();
 sg13g2_fill_8 FILLER_0_44_1014 ();
 sg13g2_fill_8 FILLER_0_44_1022 ();
 sg13g2_fill_2 FILLER_0_44_1037 ();
 sg13g2_fill_8 FILLER_0_44_1046 ();
 sg13g2_fill_8 FILLER_0_44_1054 ();
 sg13g2_fill_8 FILLER_0_44_1062 ();
 sg13g2_fill_8 FILLER_0_44_1070 ();
 sg13g2_fill_2 FILLER_0_44_1078 ();
 sg13g2_fill_1 FILLER_0_44_1080 ();
 sg13g2_fill_2 FILLER_0_44_1086 ();
 sg13g2_fill_4 FILLER_0_44_1096 ();
 sg13g2_fill_2 FILLER_0_44_1100 ();
 sg13g2_fill_1 FILLER_0_44_1102 ();
 sg13g2_fill_2 FILLER_0_44_1106 ();
 sg13g2_fill_4 FILLER_0_44_1115 ();
 sg13g2_fill_8 FILLER_0_44_1127 ();
 sg13g2_fill_8 FILLER_0_44_1135 ();
 sg13g2_fill_8 FILLER_0_44_1143 ();
 sg13g2_fill_4 FILLER_0_44_1151 ();
 sg13g2_fill_2 FILLER_0_44_1155 ();
 sg13g2_fill_8 FILLER_0_44_1163 ();
 sg13g2_fill_2 FILLER_0_44_1171 ();
 sg13g2_fill_2 FILLER_0_44_1180 ();
 sg13g2_fill_2 FILLER_0_44_1186 ();
 sg13g2_fill_2 FILLER_0_44_1193 ();
 sg13g2_fill_8 FILLER_0_44_1203 ();
 sg13g2_fill_2 FILLER_0_44_1211 ();
 sg13g2_fill_4 FILLER_0_44_1218 ();
 sg13g2_fill_2 FILLER_0_44_1222 ();
 sg13g2_fill_1 FILLER_0_44_1224 ();
 sg13g2_fill_8 FILLER_0_44_1229 ();
 sg13g2_fill_8 FILLER_0_44_1237 ();
 sg13g2_fill_8 FILLER_0_44_1245 ();
 sg13g2_fill_4 FILLER_0_44_1257 ();
 sg13g2_fill_2 FILLER_0_44_1261 ();
 sg13g2_fill_1 FILLER_0_44_1263 ();
 sg13g2_fill_4 FILLER_0_44_1269 ();
 sg13g2_fill_2 FILLER_0_44_1273 ();
 sg13g2_fill_1 FILLER_0_44_1275 ();
 sg13g2_fill_2 FILLER_0_44_1281 ();
 sg13g2_fill_4 FILLER_0_44_1288 ();
 sg13g2_fill_1 FILLER_0_44_1296 ();
 sg13g2_fill_8 FILLER_0_45_0 ();
 sg13g2_fill_8 FILLER_0_45_8 ();
 sg13g2_fill_8 FILLER_0_45_16 ();
 sg13g2_fill_8 FILLER_0_45_24 ();
 sg13g2_fill_8 FILLER_0_45_32 ();
 sg13g2_fill_8 FILLER_0_45_40 ();
 sg13g2_fill_8 FILLER_0_45_48 ();
 sg13g2_fill_8 FILLER_0_45_56 ();
 sg13g2_fill_8 FILLER_0_45_64 ();
 sg13g2_fill_8 FILLER_0_45_72 ();
 sg13g2_fill_8 FILLER_0_45_80 ();
 sg13g2_fill_8 FILLER_0_45_88 ();
 sg13g2_fill_8 FILLER_0_45_96 ();
 sg13g2_fill_8 FILLER_0_45_104 ();
 sg13g2_fill_8 FILLER_0_45_112 ();
 sg13g2_fill_8 FILLER_0_45_120 ();
 sg13g2_fill_8 FILLER_0_45_128 ();
 sg13g2_fill_8 FILLER_0_45_136 ();
 sg13g2_fill_8 FILLER_0_45_144 ();
 sg13g2_fill_8 FILLER_0_45_152 ();
 sg13g2_fill_8 FILLER_0_45_160 ();
 sg13g2_fill_8 FILLER_0_45_168 ();
 sg13g2_fill_8 FILLER_0_45_176 ();
 sg13g2_fill_8 FILLER_0_45_184 ();
 sg13g2_fill_8 FILLER_0_45_192 ();
 sg13g2_fill_8 FILLER_0_45_200 ();
 sg13g2_fill_4 FILLER_0_45_208 ();
 sg13g2_fill_8 FILLER_0_45_238 ();
 sg13g2_fill_8 FILLER_0_45_246 ();
 sg13g2_fill_8 FILLER_0_45_254 ();
 sg13g2_fill_8 FILLER_0_45_262 ();
 sg13g2_fill_8 FILLER_0_45_270 ();
 sg13g2_fill_8 FILLER_0_45_278 ();
 sg13g2_fill_8 FILLER_0_45_286 ();
 sg13g2_fill_8 FILLER_0_45_294 ();
 sg13g2_fill_8 FILLER_0_45_306 ();
 sg13g2_fill_8 FILLER_0_45_314 ();
 sg13g2_fill_8 FILLER_0_45_322 ();
 sg13g2_fill_8 FILLER_0_45_330 ();
 sg13g2_fill_8 FILLER_0_45_338 ();
 sg13g2_fill_4 FILLER_0_45_346 ();
 sg13g2_fill_2 FILLER_0_45_355 ();
 sg13g2_fill_2 FILLER_0_45_383 ();
 sg13g2_fill_1 FILLER_0_45_385 ();
 sg13g2_fill_8 FILLER_0_45_391 ();
 sg13g2_fill_4 FILLER_0_45_399 ();
 sg13g2_fill_2 FILLER_0_45_408 ();
 sg13g2_fill_2 FILLER_0_45_415 ();
 sg13g2_fill_2 FILLER_0_45_443 ();
 sg13g2_fill_1 FILLER_0_45_445 ();
 sg13g2_fill_2 FILLER_0_45_451 ();
 sg13g2_fill_1 FILLER_0_45_453 ();
 sg13g2_fill_2 FILLER_0_45_459 ();
 sg13g2_fill_1 FILLER_0_45_461 ();
 sg13g2_fill_8 FILLER_0_45_467 ();
 sg13g2_fill_8 FILLER_0_45_475 ();
 sg13g2_fill_8 FILLER_0_45_483 ();
 sg13g2_fill_8 FILLER_0_45_491 ();
 sg13g2_fill_8 FILLER_0_45_499 ();
 sg13g2_fill_2 FILLER_0_45_507 ();
 sg13g2_fill_1 FILLER_0_45_509 ();
 sg13g2_fill_2 FILLER_0_45_515 ();
 sg13g2_fill_2 FILLER_0_45_521 ();
 sg13g2_fill_8 FILLER_0_45_549 ();
 sg13g2_fill_8 FILLER_0_45_557 ();
 sg13g2_fill_8 FILLER_0_45_565 ();
 sg13g2_fill_8 FILLER_0_45_573 ();
 sg13g2_fill_8 FILLER_0_45_581 ();
 sg13g2_fill_8 FILLER_0_45_589 ();
 sg13g2_fill_8 FILLER_0_45_597 ();
 sg13g2_fill_8 FILLER_0_45_605 ();
 sg13g2_fill_8 FILLER_0_45_613 ();
 sg13g2_fill_4 FILLER_0_45_621 ();
 sg13g2_fill_1 FILLER_0_45_625 ();
 sg13g2_fill_8 FILLER_0_45_630 ();
 sg13g2_fill_8 FILLER_0_45_638 ();
 sg13g2_fill_8 FILLER_0_45_646 ();
 sg13g2_fill_8 FILLER_0_45_654 ();
 sg13g2_fill_4 FILLER_0_45_662 ();
 sg13g2_fill_2 FILLER_0_45_666 ();
 sg13g2_fill_2 FILLER_0_45_672 ();
 sg13g2_fill_8 FILLER_0_45_700 ();
 sg13g2_fill_8 FILLER_0_45_708 ();
 sg13g2_fill_4 FILLER_0_45_716 ();
 sg13g2_fill_2 FILLER_0_45_720 ();
 sg13g2_fill_8 FILLER_0_45_732 ();
 sg13g2_fill_4 FILLER_0_45_740 ();
 sg13g2_fill_2 FILLER_0_45_744 ();
 sg13g2_fill_1 FILLER_0_45_746 ();
 sg13g2_fill_8 FILLER_0_45_752 ();
 sg13g2_fill_2 FILLER_0_45_764 ();
 sg13g2_fill_2 FILLER_0_45_771 ();
 sg13g2_fill_2 FILLER_0_45_779 ();
 sg13g2_fill_4 FILLER_0_45_790 ();
 sg13g2_fill_2 FILLER_0_45_820 ();
 sg13g2_fill_4 FILLER_0_45_848 ();
 sg13g2_fill_2 FILLER_0_45_852 ();
 sg13g2_fill_4 FILLER_0_45_858 ();
 sg13g2_fill_2 FILLER_0_45_862 ();
 sg13g2_fill_4 FILLER_0_45_869 ();
 sg13g2_fill_2 FILLER_0_45_873 ();
 sg13g2_fill_8 FILLER_0_45_896 ();
 sg13g2_fill_8 FILLER_0_45_904 ();
 sg13g2_fill_8 FILLER_0_45_912 ();
 sg13g2_fill_8 FILLER_0_45_920 ();
 sg13g2_fill_8 FILLER_0_45_928 ();
 sg13g2_fill_8 FILLER_0_45_936 ();
 sg13g2_fill_8 FILLER_0_45_944 ();
 sg13g2_fill_4 FILLER_0_45_952 ();
 sg13g2_fill_2 FILLER_0_45_956 ();
 sg13g2_fill_1 FILLER_0_45_958 ();
 sg13g2_fill_2 FILLER_0_45_963 ();
 sg13g2_fill_4 FILLER_0_45_970 ();
 sg13g2_fill_2 FILLER_0_45_980 ();
 sg13g2_fill_1 FILLER_0_45_982 ();
 sg13g2_fill_2 FILLER_0_45_988 ();
 sg13g2_fill_2 FILLER_0_45_995 ();
 sg13g2_fill_2 FILLER_0_45_1002 ();
 sg13g2_fill_8 FILLER_0_45_1009 ();
 sg13g2_fill_4 FILLER_0_45_1017 ();
 sg13g2_fill_1 FILLER_0_45_1021 ();
 sg13g2_fill_2 FILLER_0_45_1027 ();
 sg13g2_fill_2 FILLER_0_45_1033 ();
 sg13g2_fill_8 FILLER_0_45_1039 ();
 sg13g2_fill_8 FILLER_0_45_1047 ();
 sg13g2_fill_8 FILLER_0_45_1055 ();
 sg13g2_fill_8 FILLER_0_45_1063 ();
 sg13g2_fill_4 FILLER_0_45_1071 ();
 sg13g2_fill_2 FILLER_0_45_1075 ();
 sg13g2_fill_1 FILLER_0_45_1077 ();
 sg13g2_fill_2 FILLER_0_45_1084 ();
 sg13g2_fill_1 FILLER_0_45_1086 ();
 sg13g2_fill_4 FILLER_0_45_1094 ();
 sg13g2_fill_2 FILLER_0_45_1098 ();
 sg13g2_fill_4 FILLER_0_45_1105 ();
 sg13g2_fill_2 FILLER_0_45_1109 ();
 sg13g2_fill_2 FILLER_0_45_1116 ();
 sg13g2_fill_2 FILLER_0_45_1123 ();
 sg13g2_fill_8 FILLER_0_45_1130 ();
 sg13g2_fill_8 FILLER_0_45_1138 ();
 sg13g2_fill_8 FILLER_0_45_1150 ();
 sg13g2_fill_8 FILLER_0_45_1163 ();
 sg13g2_fill_4 FILLER_0_45_1171 ();
 sg13g2_fill_2 FILLER_0_45_1175 ();
 sg13g2_fill_2 FILLER_0_45_1185 ();
 sg13g2_fill_2 FILLER_0_45_1195 ();
 sg13g2_fill_2 FILLER_0_45_1202 ();
 sg13g2_fill_8 FILLER_0_45_1208 ();
 sg13g2_fill_8 FILLER_0_45_1216 ();
 sg13g2_fill_8 FILLER_0_45_1224 ();
 sg13g2_fill_8 FILLER_0_45_1232 ();
 sg13g2_fill_1 FILLER_0_45_1240 ();
 sg13g2_fill_2 FILLER_0_45_1245 ();
 sg13g2_fill_1 FILLER_0_45_1247 ();
 sg13g2_fill_2 FILLER_0_45_1254 ();
 sg13g2_fill_2 FILLER_0_45_1260 ();
 sg13g2_fill_1 FILLER_0_45_1262 ();
 sg13g2_fill_2 FILLER_0_45_1268 ();
 sg13g2_fill_2 FILLER_0_45_1274 ();
 sg13g2_fill_2 FILLER_0_45_1279 ();
 sg13g2_fill_1 FILLER_0_45_1281 ();
 sg13g2_fill_4 FILLER_0_45_1287 ();
 sg13g2_fill_2 FILLER_0_45_1295 ();
 sg13g2_fill_8 FILLER_0_46_0 ();
 sg13g2_fill_8 FILLER_0_46_8 ();
 sg13g2_fill_8 FILLER_0_46_16 ();
 sg13g2_fill_8 FILLER_0_46_24 ();
 sg13g2_fill_8 FILLER_0_46_32 ();
 sg13g2_fill_8 FILLER_0_46_40 ();
 sg13g2_fill_8 FILLER_0_46_48 ();
 sg13g2_fill_8 FILLER_0_46_56 ();
 sg13g2_fill_8 FILLER_0_46_64 ();
 sg13g2_fill_8 FILLER_0_46_72 ();
 sg13g2_fill_8 FILLER_0_46_80 ();
 sg13g2_fill_8 FILLER_0_46_88 ();
 sg13g2_fill_8 FILLER_0_46_96 ();
 sg13g2_fill_8 FILLER_0_46_104 ();
 sg13g2_fill_8 FILLER_0_46_112 ();
 sg13g2_fill_8 FILLER_0_46_120 ();
 sg13g2_fill_8 FILLER_0_46_128 ();
 sg13g2_fill_8 FILLER_0_46_136 ();
 sg13g2_fill_8 FILLER_0_46_144 ();
 sg13g2_fill_8 FILLER_0_46_152 ();
 sg13g2_fill_8 FILLER_0_46_160 ();
 sg13g2_fill_8 FILLER_0_46_168 ();
 sg13g2_fill_8 FILLER_0_46_176 ();
 sg13g2_fill_8 FILLER_0_46_184 ();
 sg13g2_fill_8 FILLER_0_46_192 ();
 sg13g2_fill_8 FILLER_0_46_200 ();
 sg13g2_fill_2 FILLER_0_46_208 ();
 sg13g2_fill_8 FILLER_0_46_215 ();
 sg13g2_fill_8 FILLER_0_46_223 ();
 sg13g2_fill_8 FILLER_0_46_235 ();
 sg13g2_fill_8 FILLER_0_46_243 ();
 sg13g2_fill_4 FILLER_0_46_251 ();
 sg13g2_fill_2 FILLER_0_46_255 ();
 sg13g2_fill_1 FILLER_0_46_257 ();
 sg13g2_fill_4 FILLER_0_46_262 ();
 sg13g2_fill_1 FILLER_0_46_266 ();
 sg13g2_fill_2 FILLER_0_46_271 ();
 sg13g2_fill_4 FILLER_0_46_299 ();
 sg13g2_fill_2 FILLER_0_46_308 ();
 sg13g2_fill_8 FILLER_0_46_336 ();
 sg13g2_fill_8 FILLER_0_46_344 ();
 sg13g2_fill_2 FILLER_0_46_357 ();
 sg13g2_fill_4 FILLER_0_46_363 ();
 sg13g2_fill_8 FILLER_0_46_393 ();
 sg13g2_fill_2 FILLER_0_46_427 ();
 sg13g2_fill_2 FILLER_0_46_434 ();
 sg13g2_fill_1 FILLER_0_46_436 ();
 sg13g2_fill_2 FILLER_0_46_443 ();
 sg13g2_fill_2 FILLER_0_46_471 ();
 sg13g2_fill_4 FILLER_0_46_478 ();
 sg13g2_fill_2 FILLER_0_46_487 ();
 sg13g2_fill_2 FILLER_0_46_494 ();
 sg13g2_fill_2 FILLER_0_46_501 ();
 sg13g2_fill_2 FILLER_0_46_507 ();
 sg13g2_fill_8 FILLER_0_46_530 ();
 sg13g2_fill_8 FILLER_0_46_538 ();
 sg13g2_fill_8 FILLER_0_46_546 ();
 sg13g2_fill_8 FILLER_0_46_554 ();
 sg13g2_fill_8 FILLER_0_46_562 ();
 sg13g2_fill_4 FILLER_0_46_570 ();
 sg13g2_fill_1 FILLER_0_46_574 ();
 sg13g2_fill_8 FILLER_0_46_601 ();
 sg13g2_fill_8 FILLER_0_46_609 ();
 sg13g2_fill_4 FILLER_0_46_617 ();
 sg13g2_fill_2 FILLER_0_46_626 ();
 sg13g2_fill_2 FILLER_0_46_654 ();
 sg13g2_fill_8 FILLER_0_46_677 ();
 sg13g2_fill_8 FILLER_0_46_685 ();
 sg13g2_fill_8 FILLER_0_46_693 ();
 sg13g2_fill_8 FILLER_0_46_701 ();
 sg13g2_fill_8 FILLER_0_46_709 ();
 sg13g2_fill_8 FILLER_0_46_717 ();
 sg13g2_fill_8 FILLER_0_46_725 ();
 sg13g2_fill_2 FILLER_0_46_738 ();
 sg13g2_fill_4 FILLER_0_46_745 ();
 sg13g2_fill_1 FILLER_0_46_749 ();
 sg13g2_fill_8 FILLER_0_46_756 ();
 sg13g2_fill_8 FILLER_0_46_764 ();
 sg13g2_fill_8 FILLER_0_46_772 ();
 sg13g2_fill_8 FILLER_0_46_780 ();
 sg13g2_fill_2 FILLER_0_46_788 ();
 sg13g2_fill_1 FILLER_0_46_790 ();
 sg13g2_fill_8 FILLER_0_46_796 ();
 sg13g2_fill_4 FILLER_0_46_804 ();
 sg13g2_fill_8 FILLER_0_46_813 ();
 sg13g2_fill_2 FILLER_0_46_842 ();
 sg13g2_fill_8 FILLER_0_46_849 ();
 sg13g2_fill_2 FILLER_0_46_857 ();
 sg13g2_fill_8 FILLER_0_46_864 ();
 sg13g2_fill_4 FILLER_0_46_872 ();
 sg13g2_fill_2 FILLER_0_46_880 ();
 sg13g2_fill_2 FILLER_0_46_908 ();
 sg13g2_fill_8 FILLER_0_46_914 ();
 sg13g2_fill_8 FILLER_0_46_922 ();
 sg13g2_fill_8 FILLER_0_46_930 ();
 sg13g2_fill_8 FILLER_0_46_938 ();
 sg13g2_fill_2 FILLER_0_46_946 ();
 sg13g2_fill_2 FILLER_0_46_953 ();
 sg13g2_fill_4 FILLER_0_46_961 ();
 sg13g2_fill_2 FILLER_0_46_965 ();
 sg13g2_fill_2 FILLER_0_46_972 ();
 sg13g2_fill_1 FILLER_0_46_974 ();
 sg13g2_fill_8 FILLER_0_46_980 ();
 sg13g2_fill_2 FILLER_0_46_988 ();
 sg13g2_fill_2 FILLER_0_46_995 ();
 sg13g2_fill_2 FILLER_0_46_1001 ();
 sg13g2_fill_1 FILLER_0_46_1003 ();
 sg13g2_fill_8 FILLER_0_46_1009 ();
 sg13g2_fill_8 FILLER_0_46_1017 ();
 sg13g2_fill_1 FILLER_0_46_1025 ();
 sg13g2_fill_2 FILLER_0_46_1032 ();
 sg13g2_fill_2 FILLER_0_46_1040 ();
 sg13g2_fill_8 FILLER_0_46_1045 ();
 sg13g2_fill_8 FILLER_0_46_1053 ();
 sg13g2_fill_8 FILLER_0_46_1061 ();
 sg13g2_fill_2 FILLER_0_46_1069 ();
 sg13g2_fill_1 FILLER_0_46_1071 ();
 sg13g2_fill_8 FILLER_0_46_1077 ();
 sg13g2_fill_4 FILLER_0_46_1085 ();
 sg13g2_fill_2 FILLER_0_46_1089 ();
 sg13g2_fill_2 FILLER_0_46_1096 ();
 sg13g2_fill_2 FILLER_0_46_1102 ();
 sg13g2_fill_2 FILLER_0_46_1112 ();
 sg13g2_fill_4 FILLER_0_46_1117 ();
 sg13g2_fill_2 FILLER_0_46_1121 ();
 sg13g2_fill_2 FILLER_0_46_1129 ();
 sg13g2_fill_1 FILLER_0_46_1131 ();
 sg13g2_fill_2 FILLER_0_46_1136 ();
 sg13g2_fill_2 FILLER_0_46_1143 ();
 sg13g2_fill_1 FILLER_0_46_1145 ();
 sg13g2_fill_4 FILLER_0_46_1151 ();
 sg13g2_fill_8 FILLER_0_46_1161 ();
 sg13g2_fill_8 FILLER_0_46_1169 ();
 sg13g2_fill_1 FILLER_0_46_1177 ();
 sg13g2_fill_8 FILLER_0_46_1182 ();
 sg13g2_fill_2 FILLER_0_46_1190 ();
 sg13g2_fill_1 FILLER_0_46_1192 ();
 sg13g2_fill_4 FILLER_0_46_1198 ();
 sg13g2_fill_2 FILLER_0_46_1202 ();
 sg13g2_fill_4 FILLER_0_46_1212 ();
 sg13g2_fill_2 FILLER_0_46_1216 ();
 sg13g2_fill_2 FILLER_0_46_1224 ();
 sg13g2_fill_8 FILLER_0_46_1231 ();
 sg13g2_fill_4 FILLER_0_46_1239 ();
 sg13g2_fill_8 FILLER_0_46_1248 ();
 sg13g2_fill_2 FILLER_0_46_1261 ();
 sg13g2_fill_4 FILLER_0_46_1268 ();
 sg13g2_fill_8 FILLER_0_46_1277 ();
 sg13g2_fill_1 FILLER_0_46_1285 ();
 sg13g2_fill_2 FILLER_0_46_1290 ();
 sg13g2_fill_1 FILLER_0_46_1296 ();
 sg13g2_fill_8 FILLER_0_47_0 ();
 sg13g2_fill_8 FILLER_0_47_8 ();
 sg13g2_fill_8 FILLER_0_47_16 ();
 sg13g2_fill_8 FILLER_0_47_24 ();
 sg13g2_fill_8 FILLER_0_47_32 ();
 sg13g2_fill_8 FILLER_0_47_40 ();
 sg13g2_fill_8 FILLER_0_47_48 ();
 sg13g2_fill_8 FILLER_0_47_56 ();
 sg13g2_fill_8 FILLER_0_47_64 ();
 sg13g2_fill_8 FILLER_0_47_72 ();
 sg13g2_fill_8 FILLER_0_47_80 ();
 sg13g2_fill_8 FILLER_0_47_88 ();
 sg13g2_fill_8 FILLER_0_47_96 ();
 sg13g2_fill_8 FILLER_0_47_104 ();
 sg13g2_fill_8 FILLER_0_47_112 ();
 sg13g2_fill_8 FILLER_0_47_120 ();
 sg13g2_fill_8 FILLER_0_47_128 ();
 sg13g2_fill_8 FILLER_0_47_136 ();
 sg13g2_fill_8 FILLER_0_47_144 ();
 sg13g2_fill_8 FILLER_0_47_152 ();
 sg13g2_fill_8 FILLER_0_47_160 ();
 sg13g2_fill_8 FILLER_0_47_168 ();
 sg13g2_fill_8 FILLER_0_47_176 ();
 sg13g2_fill_8 FILLER_0_47_184 ();
 sg13g2_fill_8 FILLER_0_47_192 ();
 sg13g2_fill_8 FILLER_0_47_200 ();
 sg13g2_fill_8 FILLER_0_47_208 ();
 sg13g2_fill_8 FILLER_0_47_216 ();
 sg13g2_fill_8 FILLER_0_47_224 ();
 sg13g2_fill_8 FILLER_0_47_232 ();
 sg13g2_fill_8 FILLER_0_47_240 ();
 sg13g2_fill_4 FILLER_0_47_253 ();
 sg13g2_fill_2 FILLER_0_47_262 ();
 sg13g2_fill_2 FILLER_0_47_269 ();
 sg13g2_fill_2 FILLER_0_47_297 ();
 sg13g2_fill_2 FILLER_0_47_309 ();
 sg13g2_fill_2 FILLER_0_47_315 ();
 sg13g2_fill_8 FILLER_0_47_343 ();
 sg13g2_fill_1 FILLER_0_47_351 ();
 sg13g2_fill_8 FILLER_0_47_357 ();
 sg13g2_fill_4 FILLER_0_47_365 ();
 sg13g2_fill_2 FILLER_0_47_369 ();
 sg13g2_fill_1 FILLER_0_47_371 ();
 sg13g2_fill_2 FILLER_0_47_377 ();
 sg13g2_fill_8 FILLER_0_47_389 ();
 sg13g2_fill_8 FILLER_0_47_397 ();
 sg13g2_fill_4 FILLER_0_47_405 ();
 sg13g2_fill_4 FILLER_0_47_413 ();
 sg13g2_fill_8 FILLER_0_47_422 ();
 sg13g2_fill_8 FILLER_0_47_430 ();
 sg13g2_fill_8 FILLER_0_47_438 ();
 sg13g2_fill_8 FILLER_0_47_446 ();
 sg13g2_fill_2 FILLER_0_47_454 ();
 sg13g2_fill_8 FILLER_0_47_461 ();
 sg13g2_fill_2 FILLER_0_47_469 ();
 sg13g2_fill_1 FILLER_0_47_471 ();
 sg13g2_fill_8 FILLER_0_47_479 ();
 sg13g2_fill_1 FILLER_0_47_487 ();
 sg13g2_fill_2 FILLER_0_47_493 ();
 sg13g2_fill_4 FILLER_0_47_500 ();
 sg13g2_fill_8 FILLER_0_47_530 ();
 sg13g2_fill_8 FILLER_0_47_538 ();
 sg13g2_fill_8 FILLER_0_47_546 ();
 sg13g2_fill_8 FILLER_0_47_554 ();
 sg13g2_fill_8 FILLER_0_47_562 ();
 sg13g2_fill_2 FILLER_0_47_575 ();
 sg13g2_fill_2 FILLER_0_47_581 ();
 sg13g2_fill_1 FILLER_0_47_583 ();
 sg13g2_fill_4 FILLER_0_47_589 ();
 sg13g2_fill_2 FILLER_0_47_593 ();
 sg13g2_fill_1 FILLER_0_47_595 ();
 sg13g2_fill_2 FILLER_0_47_600 ();
 sg13g2_fill_2 FILLER_0_47_623 ();
 sg13g2_fill_8 FILLER_0_47_629 ();
 sg13g2_fill_4 FILLER_0_47_637 ();
 sg13g2_fill_1 FILLER_0_47_641 ();
 sg13g2_fill_2 FILLER_0_47_647 ();
 sg13g2_fill_2 FILLER_0_47_653 ();
 sg13g2_fill_1 FILLER_0_47_655 ();
 sg13g2_fill_8 FILLER_0_47_677 ();
 sg13g2_fill_4 FILLER_0_47_685 ();
 sg13g2_fill_4 FILLER_0_47_694 ();
 sg13g2_fill_1 FILLER_0_47_698 ();
 sg13g2_fill_4 FILLER_0_47_703 ();
 sg13g2_fill_1 FILLER_0_47_707 ();
 sg13g2_fill_4 FILLER_0_47_713 ();
 sg13g2_fill_2 FILLER_0_47_717 ();
 sg13g2_fill_8 FILLER_0_47_724 ();
 sg13g2_fill_1 FILLER_0_47_732 ();
 sg13g2_fill_8 FILLER_0_47_743 ();
 sg13g2_fill_8 FILLER_0_47_751 ();
 sg13g2_fill_4 FILLER_0_47_759 ();
 sg13g2_fill_2 FILLER_0_47_771 ();
 sg13g2_fill_8 FILLER_0_47_778 ();
 sg13g2_fill_8 FILLER_0_47_786 ();
 sg13g2_fill_4 FILLER_0_47_794 ();
 sg13g2_fill_1 FILLER_0_47_798 ();
 sg13g2_fill_2 FILLER_0_47_825 ();
 sg13g2_fill_8 FILLER_0_47_832 ();
 sg13g2_fill_8 FILLER_0_47_840 ();
 sg13g2_fill_8 FILLER_0_47_848 ();
 sg13g2_fill_2 FILLER_0_47_856 ();
 sg13g2_fill_2 FILLER_0_47_884 ();
 sg13g2_fill_2 FILLER_0_47_907 ();
 sg13g2_fill_8 FILLER_0_47_914 ();
 sg13g2_fill_8 FILLER_0_47_922 ();
 sg13g2_fill_8 FILLER_0_47_930 ();
 sg13g2_fill_4 FILLER_0_47_942 ();
 sg13g2_fill_1 FILLER_0_47_946 ();
 sg13g2_fill_2 FILLER_0_47_953 ();
 sg13g2_fill_2 FILLER_0_47_961 ();
 sg13g2_fill_8 FILLER_0_47_968 ();
 sg13g2_fill_8 FILLER_0_47_976 ();
 sg13g2_fill_8 FILLER_0_47_984 ();
 sg13g2_fill_2 FILLER_0_47_992 ();
 sg13g2_fill_2 FILLER_0_47_999 ();
 sg13g2_fill_1 FILLER_0_47_1001 ();
 sg13g2_fill_8 FILLER_0_47_1009 ();
 sg13g2_fill_4 FILLER_0_47_1017 ();
 sg13g2_fill_2 FILLER_0_47_1021 ();
 sg13g2_fill_2 FILLER_0_47_1028 ();
 sg13g2_fill_8 FILLER_0_47_1035 ();
 sg13g2_fill_8 FILLER_0_47_1043 ();
 sg13g2_fill_8 FILLER_0_47_1051 ();
 sg13g2_fill_8 FILLER_0_47_1059 ();
 sg13g2_fill_4 FILLER_0_47_1067 ();
 sg13g2_fill_1 FILLER_0_47_1071 ();
 sg13g2_fill_8 FILLER_0_47_1082 ();
 sg13g2_fill_4 FILLER_0_47_1090 ();
 sg13g2_fill_2 FILLER_0_47_1099 ();
 sg13g2_fill_4 FILLER_0_47_1105 ();
 sg13g2_fill_2 FILLER_0_47_1109 ();
 sg13g2_fill_2 FILLER_0_47_1118 ();
 sg13g2_fill_8 FILLER_0_47_1125 ();
 sg13g2_fill_4 FILLER_0_47_1133 ();
 sg13g2_fill_2 FILLER_0_47_1137 ();
 sg13g2_fill_8 FILLER_0_47_1147 ();
 sg13g2_fill_1 FILLER_0_47_1155 ();
 sg13g2_fill_8 FILLER_0_47_1161 ();
 sg13g2_fill_4 FILLER_0_47_1169 ();
 sg13g2_fill_4 FILLER_0_47_1178 ();
 sg13g2_fill_2 FILLER_0_47_1187 ();
 sg13g2_fill_1 FILLER_0_47_1189 ();
 sg13g2_fill_2 FILLER_0_47_1198 ();
 sg13g2_fill_4 FILLER_0_47_1203 ();
 sg13g2_fill_2 FILLER_0_47_1207 ();
 sg13g2_fill_1 FILLER_0_47_1209 ();
 sg13g2_fill_2 FILLER_0_47_1215 ();
 sg13g2_fill_8 FILLER_0_47_1221 ();
 sg13g2_fill_8 FILLER_0_47_1229 ();
 sg13g2_fill_8 FILLER_0_47_1245 ();
 sg13g2_fill_2 FILLER_0_47_1257 ();
 sg13g2_fill_8 FILLER_0_47_1263 ();
 sg13g2_fill_4 FILLER_0_47_1271 ();
 sg13g2_fill_2 FILLER_0_47_1275 ();
 sg13g2_fill_8 FILLER_0_47_1281 ();
 sg13g2_fill_2 FILLER_0_47_1289 ();
 sg13g2_fill_2 FILLER_0_47_1295 ();
 sg13g2_fill_8 FILLER_0_48_0 ();
 sg13g2_fill_8 FILLER_0_48_8 ();
 sg13g2_fill_8 FILLER_0_48_16 ();
 sg13g2_fill_8 FILLER_0_48_24 ();
 sg13g2_fill_8 FILLER_0_48_32 ();
 sg13g2_fill_8 FILLER_0_48_40 ();
 sg13g2_fill_8 FILLER_0_48_48 ();
 sg13g2_fill_8 FILLER_0_48_56 ();
 sg13g2_fill_8 FILLER_0_48_64 ();
 sg13g2_fill_8 FILLER_0_48_72 ();
 sg13g2_fill_8 FILLER_0_48_80 ();
 sg13g2_fill_8 FILLER_0_48_88 ();
 sg13g2_fill_8 FILLER_0_48_96 ();
 sg13g2_fill_8 FILLER_0_48_104 ();
 sg13g2_fill_8 FILLER_0_48_112 ();
 sg13g2_fill_8 FILLER_0_48_120 ();
 sg13g2_fill_8 FILLER_0_48_128 ();
 sg13g2_fill_8 FILLER_0_48_136 ();
 sg13g2_fill_8 FILLER_0_48_144 ();
 sg13g2_fill_8 FILLER_0_48_152 ();
 sg13g2_fill_8 FILLER_0_48_160 ();
 sg13g2_fill_8 FILLER_0_48_168 ();
 sg13g2_fill_8 FILLER_0_48_176 ();
 sg13g2_fill_8 FILLER_0_48_184 ();
 sg13g2_fill_8 FILLER_0_48_192 ();
 sg13g2_fill_8 FILLER_0_48_200 ();
 sg13g2_fill_8 FILLER_0_48_208 ();
 sg13g2_fill_8 FILLER_0_48_216 ();
 sg13g2_fill_8 FILLER_0_48_224 ();
 sg13g2_fill_8 FILLER_0_48_232 ();
 sg13g2_fill_1 FILLER_0_48_240 ();
 sg13g2_fill_4 FILLER_0_48_267 ();
 sg13g2_fill_2 FILLER_0_48_271 ();
 sg13g2_fill_4 FILLER_0_48_278 ();
 sg13g2_fill_1 FILLER_0_48_282 ();
 sg13g2_fill_4 FILLER_0_48_288 ();
 sg13g2_fill_2 FILLER_0_48_313 ();
 sg13g2_fill_1 FILLER_0_48_315 ();
 sg13g2_fill_4 FILLER_0_48_321 ();
 sg13g2_fill_4 FILLER_0_48_330 ();
 sg13g2_fill_2 FILLER_0_48_344 ();
 sg13g2_fill_4 FILLER_0_48_350 ();
 sg13g2_fill_2 FILLER_0_48_354 ();
 sg13g2_fill_1 FILLER_0_48_356 ();
 sg13g2_fill_2 FILLER_0_48_362 ();
 sg13g2_fill_4 FILLER_0_48_369 ();
 sg13g2_fill_8 FILLER_0_48_377 ();
 sg13g2_fill_8 FILLER_0_48_385 ();
 sg13g2_fill_2 FILLER_0_48_393 ();
 sg13g2_fill_8 FILLER_0_48_400 ();
 sg13g2_fill_4 FILLER_0_48_408 ();
 sg13g2_fill_2 FILLER_0_48_412 ();
 sg13g2_fill_4 FILLER_0_48_420 ();
 sg13g2_fill_1 FILLER_0_48_424 ();
 sg13g2_fill_8 FILLER_0_48_433 ();
 sg13g2_fill_4 FILLER_0_48_441 ();
 sg13g2_fill_1 FILLER_0_48_445 ();
 sg13g2_fill_4 FILLER_0_48_454 ();
 sg13g2_fill_4 FILLER_0_48_463 ();
 sg13g2_fill_4 FILLER_0_48_471 ();
 sg13g2_fill_8 FILLER_0_48_480 ();
 sg13g2_fill_8 FILLER_0_48_488 ();
 sg13g2_fill_8 FILLER_0_48_496 ();
 sg13g2_fill_2 FILLER_0_48_504 ();
 sg13g2_fill_8 FILLER_0_48_532 ();
 sg13g2_fill_8 FILLER_0_48_540 ();
 sg13g2_fill_8 FILLER_0_48_548 ();
 sg13g2_fill_8 FILLER_0_48_560 ();
 sg13g2_fill_2 FILLER_0_48_573 ();
 sg13g2_fill_4 FILLER_0_48_601 ();
 sg13g2_fill_1 FILLER_0_48_605 ();
 sg13g2_fill_4 FILLER_0_48_632 ();
 sg13g2_fill_2 FILLER_0_48_636 ();
 sg13g2_fill_1 FILLER_0_48_638 ();
 sg13g2_fill_2 FILLER_0_48_665 ();
 sg13g2_fill_2 FILLER_0_48_672 ();
 sg13g2_fill_2 FILLER_0_48_679 ();
 sg13g2_fill_2 FILLER_0_48_686 ();
 sg13g2_fill_4 FILLER_0_48_714 ();
 sg13g2_fill_1 FILLER_0_48_718 ();
 sg13g2_fill_2 FILLER_0_48_745 ();
 sg13g2_fill_1 FILLER_0_48_747 ();
 sg13g2_fill_2 FILLER_0_48_774 ();
 sg13g2_fill_1 FILLER_0_48_776 ();
 sg13g2_fill_8 FILLER_0_48_781 ();
 sg13g2_fill_2 FILLER_0_48_789 ();
 sg13g2_fill_1 FILLER_0_48_791 ();
 sg13g2_fill_2 FILLER_0_48_797 ();
 sg13g2_fill_2 FILLER_0_48_825 ();
 sg13g2_fill_2 FILLER_0_48_831 ();
 sg13g2_fill_8 FILLER_0_48_838 ();
 sg13g2_fill_8 FILLER_0_48_846 ();
 sg13g2_fill_2 FILLER_0_48_854 ();
 sg13g2_fill_1 FILLER_0_48_856 ();
 sg13g2_fill_2 FILLER_0_48_862 ();
 sg13g2_fill_4 FILLER_0_48_869 ();
 sg13g2_fill_4 FILLER_0_48_899 ();
 sg13g2_fill_2 FILLER_0_48_903 ();
 sg13g2_fill_1 FILLER_0_48_905 ();
 sg13g2_fill_8 FILLER_0_48_910 ();
 sg13g2_fill_8 FILLER_0_48_918 ();
 sg13g2_fill_2 FILLER_0_48_926 ();
 sg13g2_fill_1 FILLER_0_48_928 ();
 sg13g2_fill_8 FILLER_0_48_933 ();
 sg13g2_fill_4 FILLER_0_48_941 ();
 sg13g2_fill_2 FILLER_0_48_945 ();
 sg13g2_fill_2 FILLER_0_48_953 ();
 sg13g2_fill_2 FILLER_0_48_961 ();
 sg13g2_fill_8 FILLER_0_48_967 ();
 sg13g2_fill_8 FILLER_0_48_975 ();
 sg13g2_fill_8 FILLER_0_48_983 ();
 sg13g2_fill_2 FILLER_0_48_991 ();
 sg13g2_fill_2 FILLER_0_48_1001 ();
 sg13g2_fill_8 FILLER_0_48_1008 ();
 sg13g2_fill_8 FILLER_0_48_1016 ();
 sg13g2_fill_8 FILLER_0_48_1024 ();
 sg13g2_fill_2 FILLER_0_48_1032 ();
 sg13g2_fill_1 FILLER_0_48_1034 ();
 sg13g2_fill_2 FILLER_0_48_1040 ();
 sg13g2_fill_8 FILLER_0_48_1046 ();
 sg13g2_fill_8 FILLER_0_48_1054 ();
 sg13g2_fill_8 FILLER_0_48_1062 ();
 sg13g2_fill_1 FILLER_0_48_1070 ();
 sg13g2_fill_8 FILLER_0_48_1079 ();
 sg13g2_fill_1 FILLER_0_48_1087 ();
 sg13g2_fill_8 FILLER_0_48_1093 ();
 sg13g2_fill_1 FILLER_0_48_1101 ();
 sg13g2_fill_2 FILLER_0_48_1107 ();
 sg13g2_fill_2 FILLER_0_48_1114 ();
 sg13g2_fill_2 FILLER_0_48_1126 ();
 sg13g2_fill_8 FILLER_0_48_1133 ();
 sg13g2_fill_4 FILLER_0_48_1141 ();
 sg13g2_fill_1 FILLER_0_48_1145 ();
 sg13g2_fill_2 FILLER_0_48_1151 ();
 sg13g2_fill_8 FILLER_0_48_1158 ();
 sg13g2_fill_8 FILLER_0_48_1166 ();
 sg13g2_fill_1 FILLER_0_48_1174 ();
 sg13g2_fill_2 FILLER_0_48_1180 ();
 sg13g2_fill_4 FILLER_0_48_1186 ();
 sg13g2_fill_1 FILLER_0_48_1190 ();
 sg13g2_fill_2 FILLER_0_48_1199 ();
 sg13g2_fill_2 FILLER_0_48_1204 ();
 sg13g2_fill_8 FILLER_0_48_1214 ();
 sg13g2_fill_2 FILLER_0_48_1226 ();
 sg13g2_fill_1 FILLER_0_48_1228 ();
 sg13g2_fill_2 FILLER_0_48_1234 ();
 sg13g2_fill_2 FILLER_0_48_1241 ();
 sg13g2_fill_1 FILLER_0_48_1243 ();
 sg13g2_fill_8 FILLER_0_48_1249 ();
 sg13g2_fill_2 FILLER_0_48_1257 ();
 sg13g2_fill_4 FILLER_0_48_1263 ();
 sg13g2_fill_2 FILLER_0_48_1272 ();
 sg13g2_fill_2 FILLER_0_48_1279 ();
 sg13g2_fill_8 FILLER_0_48_1286 ();
 sg13g2_fill_2 FILLER_0_48_1294 ();
 sg13g2_fill_1 FILLER_0_48_1296 ();
 sg13g2_fill_8 FILLER_0_49_0 ();
 sg13g2_fill_8 FILLER_0_49_8 ();
 sg13g2_fill_8 FILLER_0_49_16 ();
 sg13g2_fill_8 FILLER_0_49_24 ();
 sg13g2_fill_8 FILLER_0_49_32 ();
 sg13g2_fill_8 FILLER_0_49_40 ();
 sg13g2_fill_8 FILLER_0_49_48 ();
 sg13g2_fill_8 FILLER_0_49_56 ();
 sg13g2_fill_8 FILLER_0_49_64 ();
 sg13g2_fill_8 FILLER_0_49_72 ();
 sg13g2_fill_8 FILLER_0_49_80 ();
 sg13g2_fill_8 FILLER_0_49_88 ();
 sg13g2_fill_8 FILLER_0_49_96 ();
 sg13g2_fill_8 FILLER_0_49_104 ();
 sg13g2_fill_8 FILLER_0_49_112 ();
 sg13g2_fill_8 FILLER_0_49_120 ();
 sg13g2_fill_8 FILLER_0_49_128 ();
 sg13g2_fill_8 FILLER_0_49_136 ();
 sg13g2_fill_8 FILLER_0_49_144 ();
 sg13g2_fill_8 FILLER_0_49_152 ();
 sg13g2_fill_8 FILLER_0_49_160 ();
 sg13g2_fill_8 FILLER_0_49_168 ();
 sg13g2_fill_8 FILLER_0_49_176 ();
 sg13g2_fill_8 FILLER_0_49_184 ();
 sg13g2_fill_8 FILLER_0_49_192 ();
 sg13g2_fill_8 FILLER_0_49_200 ();
 sg13g2_fill_8 FILLER_0_49_208 ();
 sg13g2_fill_8 FILLER_0_49_216 ();
 sg13g2_fill_1 FILLER_0_49_224 ();
 sg13g2_fill_2 FILLER_0_49_230 ();
 sg13g2_fill_8 FILLER_0_49_236 ();
 sg13g2_fill_2 FILLER_0_49_244 ();
 sg13g2_fill_1 FILLER_0_49_246 ();
 sg13g2_fill_2 FILLER_0_49_251 ();
 sg13g2_fill_8 FILLER_0_49_258 ();
 sg13g2_fill_4 FILLER_0_49_266 ();
 sg13g2_fill_2 FILLER_0_49_275 ();
 sg13g2_fill_2 FILLER_0_49_282 ();
 sg13g2_fill_8 FILLER_0_49_288 ();
 sg13g2_fill_8 FILLER_0_49_296 ();
 sg13g2_fill_8 FILLER_0_49_304 ();
 sg13g2_fill_2 FILLER_0_49_312 ();
 sg13g2_fill_8 FILLER_0_49_319 ();
 sg13g2_fill_8 FILLER_0_49_327 ();
 sg13g2_fill_8 FILLER_0_49_335 ();
 sg13g2_fill_8 FILLER_0_49_343 ();
 sg13g2_fill_8 FILLER_0_49_351 ();
 sg13g2_fill_2 FILLER_0_49_359 ();
 sg13g2_fill_8 FILLER_0_49_367 ();
 sg13g2_fill_1 FILLER_0_49_375 ();
 sg13g2_fill_2 FILLER_0_49_386 ();
 sg13g2_fill_8 FILLER_0_49_394 ();
 sg13g2_fill_4 FILLER_0_49_407 ();
 sg13g2_fill_2 FILLER_0_49_411 ();
 sg13g2_fill_1 FILLER_0_49_413 ();
 sg13g2_fill_8 FILLER_0_49_420 ();
 sg13g2_fill_2 FILLER_0_49_428 ();
 sg13g2_fill_2 FILLER_0_49_436 ();
 sg13g2_fill_2 FILLER_0_49_442 ();
 sg13g2_fill_2 FILLER_0_49_470 ();
 sg13g2_fill_8 FILLER_0_49_477 ();
 sg13g2_fill_8 FILLER_0_49_485 ();
 sg13g2_fill_8 FILLER_0_49_493 ();
 sg13g2_fill_8 FILLER_0_49_501 ();
 sg13g2_fill_2 FILLER_0_49_509 ();
 sg13g2_fill_2 FILLER_0_49_516 ();
 sg13g2_fill_8 FILLER_0_49_528 ();
 sg13g2_fill_4 FILLER_0_49_536 ();
 sg13g2_fill_2 FILLER_0_49_540 ();
 sg13g2_fill_1 FILLER_0_49_542 ();
 sg13g2_fill_2 FILLER_0_49_548 ();
 sg13g2_fill_2 FILLER_0_49_555 ();
 sg13g2_fill_8 FILLER_0_49_583 ();
 sg13g2_fill_4 FILLER_0_49_591 ();
 sg13g2_fill_4 FILLER_0_49_616 ();
 sg13g2_fill_8 FILLER_0_49_625 ();
 sg13g2_fill_8 FILLER_0_49_633 ();
 sg13g2_fill_8 FILLER_0_49_641 ();
 sg13g2_fill_8 FILLER_0_49_649 ();
 sg13g2_fill_4 FILLER_0_49_657 ();
 sg13g2_fill_2 FILLER_0_49_661 ();
 sg13g2_fill_1 FILLER_0_49_663 ();
 sg13g2_fill_8 FILLER_0_49_674 ();
 sg13g2_fill_8 FILLER_0_49_682 ();
 sg13g2_fill_8 FILLER_0_49_690 ();
 sg13g2_fill_8 FILLER_0_49_698 ();
 sg13g2_fill_8 FILLER_0_49_706 ();
 sg13g2_fill_4 FILLER_0_49_714 ();
 sg13g2_fill_1 FILLER_0_49_718 ();
 sg13g2_fill_8 FILLER_0_49_723 ();
 sg13g2_fill_8 FILLER_0_49_731 ();
 sg13g2_fill_8 FILLER_0_49_739 ();
 sg13g2_fill_8 FILLER_0_49_747 ();
 sg13g2_fill_8 FILLER_0_49_755 ();
 sg13g2_fill_8 FILLER_0_49_763 ();
 sg13g2_fill_8 FILLER_0_49_771 ();
 sg13g2_fill_2 FILLER_0_49_779 ();
 sg13g2_fill_1 FILLER_0_49_781 ();
 sg13g2_fill_8 FILLER_0_49_787 ();
 sg13g2_fill_8 FILLER_0_49_799 ();
 sg13g2_fill_8 FILLER_0_49_807 ();
 sg13g2_fill_1 FILLER_0_49_815 ();
 sg13g2_fill_4 FILLER_0_49_826 ();
 sg13g2_fill_2 FILLER_0_49_830 ();
 sg13g2_fill_1 FILLER_0_49_832 ();
 sg13g2_fill_2 FILLER_0_49_838 ();
 sg13g2_fill_2 FILLER_0_49_866 ();
 sg13g2_fill_2 FILLER_0_49_872 ();
 sg13g2_fill_4 FILLER_0_49_879 ();
 sg13g2_fill_2 FILLER_0_49_883 ();
 sg13g2_fill_8 FILLER_0_49_889 ();
 sg13g2_fill_8 FILLER_0_49_897 ();
 sg13g2_fill_8 FILLER_0_49_905 ();
 sg13g2_fill_8 FILLER_0_49_913 ();
 sg13g2_fill_8 FILLER_0_49_921 ();
 sg13g2_fill_8 FILLER_0_49_929 ();
 sg13g2_fill_8 FILLER_0_49_937 ();
 sg13g2_fill_4 FILLER_0_49_945 ();
 sg13g2_fill_2 FILLER_0_49_954 ();
 sg13g2_fill_8 FILLER_0_49_960 ();
 sg13g2_fill_8 FILLER_0_49_968 ();
 sg13g2_fill_4 FILLER_0_49_976 ();
 sg13g2_fill_2 FILLER_0_49_980 ();
 sg13g2_fill_1 FILLER_0_49_982 ();
 sg13g2_fill_8 FILLER_0_49_988 ();
 sg13g2_fill_8 FILLER_0_49_996 ();
 sg13g2_fill_8 FILLER_0_49_1004 ();
 sg13g2_fill_8 FILLER_0_49_1012 ();
 sg13g2_fill_8 FILLER_0_49_1020 ();
 sg13g2_fill_8 FILLER_0_49_1028 ();
 sg13g2_fill_8 FILLER_0_49_1036 ();
 sg13g2_fill_8 FILLER_0_49_1044 ();
 sg13g2_fill_8 FILLER_0_49_1052 ();
 sg13g2_fill_8 FILLER_0_49_1060 ();
 sg13g2_fill_4 FILLER_0_49_1068 ();
 sg13g2_fill_4 FILLER_0_49_1077 ();
 sg13g2_fill_2 FILLER_0_49_1081 ();
 sg13g2_fill_8 FILLER_0_49_1089 ();
 sg13g2_fill_8 FILLER_0_49_1097 ();
 sg13g2_fill_1 FILLER_0_49_1105 ();
 sg13g2_fill_2 FILLER_0_49_1110 ();
 sg13g2_fill_8 FILLER_0_49_1118 ();
 sg13g2_fill_4 FILLER_0_49_1126 ();
 sg13g2_fill_1 FILLER_0_49_1130 ();
 sg13g2_fill_2 FILLER_0_49_1135 ();
 sg13g2_fill_2 FILLER_0_49_1142 ();
 sg13g2_fill_8 FILLER_0_49_1153 ();
 sg13g2_fill_8 FILLER_0_49_1161 ();
 sg13g2_fill_8 FILLER_0_49_1169 ();
 sg13g2_fill_2 FILLER_0_49_1177 ();
 sg13g2_fill_1 FILLER_0_49_1179 ();
 sg13g2_fill_4 FILLER_0_49_1185 ();
 sg13g2_fill_2 FILLER_0_49_1189 ();
 sg13g2_fill_4 FILLER_0_49_1199 ();
 sg13g2_fill_2 FILLER_0_49_1203 ();
 sg13g2_fill_8 FILLER_0_49_1210 ();
 sg13g2_fill_8 FILLER_0_49_1218 ();
 sg13g2_fill_8 FILLER_0_49_1226 ();
 sg13g2_fill_2 FILLER_0_49_1234 ();
 sg13g2_fill_2 FILLER_0_49_1243 ();
 sg13g2_fill_1 FILLER_0_49_1245 ();
 sg13g2_fill_2 FILLER_0_49_1251 ();
 sg13g2_fill_4 FILLER_0_49_1258 ();
 sg13g2_fill_2 FILLER_0_49_1262 ();
 sg13g2_fill_1 FILLER_0_49_1264 ();
 sg13g2_fill_8 FILLER_0_49_1269 ();
 sg13g2_fill_2 FILLER_0_49_1277 ();
 sg13g2_fill_8 FILLER_0_49_1284 ();
 sg13g2_fill_1 FILLER_0_49_1296 ();
 sg13g2_fill_8 FILLER_0_50_0 ();
 sg13g2_fill_8 FILLER_0_50_8 ();
 sg13g2_fill_8 FILLER_0_50_16 ();
 sg13g2_fill_8 FILLER_0_50_24 ();
 sg13g2_fill_8 FILLER_0_50_32 ();
 sg13g2_fill_8 FILLER_0_50_40 ();
 sg13g2_fill_8 FILLER_0_50_48 ();
 sg13g2_fill_8 FILLER_0_50_56 ();
 sg13g2_fill_8 FILLER_0_50_64 ();
 sg13g2_fill_8 FILLER_0_50_72 ();
 sg13g2_fill_8 FILLER_0_50_80 ();
 sg13g2_fill_8 FILLER_0_50_88 ();
 sg13g2_fill_8 FILLER_0_50_96 ();
 sg13g2_fill_8 FILLER_0_50_104 ();
 sg13g2_fill_8 FILLER_0_50_112 ();
 sg13g2_fill_8 FILLER_0_50_120 ();
 sg13g2_fill_8 FILLER_0_50_128 ();
 sg13g2_fill_8 FILLER_0_50_136 ();
 sg13g2_fill_8 FILLER_0_50_144 ();
 sg13g2_fill_8 FILLER_0_50_152 ();
 sg13g2_fill_8 FILLER_0_50_160 ();
 sg13g2_fill_8 FILLER_0_50_168 ();
 sg13g2_fill_8 FILLER_0_50_176 ();
 sg13g2_fill_8 FILLER_0_50_184 ();
 sg13g2_fill_8 FILLER_0_50_192 ();
 sg13g2_fill_8 FILLER_0_50_200 ();
 sg13g2_fill_8 FILLER_0_50_208 ();
 sg13g2_fill_2 FILLER_0_50_216 ();
 sg13g2_fill_1 FILLER_0_50_218 ();
 sg13g2_fill_2 FILLER_0_50_245 ();
 sg13g2_fill_1 FILLER_0_50_247 ();
 sg13g2_fill_8 FILLER_0_50_269 ();
 sg13g2_fill_8 FILLER_0_50_277 ();
 sg13g2_fill_8 FILLER_0_50_285 ();
 sg13g2_fill_8 FILLER_0_50_293 ();
 sg13g2_fill_8 FILLER_0_50_301 ();
 sg13g2_fill_8 FILLER_0_50_309 ();
 sg13g2_fill_8 FILLER_0_50_317 ();
 sg13g2_fill_8 FILLER_0_50_330 ();
 sg13g2_fill_1 FILLER_0_50_338 ();
 sg13g2_fill_2 FILLER_0_50_344 ();
 sg13g2_fill_8 FILLER_0_50_350 ();
 sg13g2_fill_4 FILLER_0_50_358 ();
 sg13g2_fill_2 FILLER_0_50_367 ();
 sg13g2_fill_8 FILLER_0_50_375 ();
 sg13g2_fill_4 FILLER_0_50_383 ();
 sg13g2_fill_8 FILLER_0_50_392 ();
 sg13g2_fill_8 FILLER_0_50_400 ();
 sg13g2_fill_8 FILLER_0_50_408 ();
 sg13g2_fill_8 FILLER_0_50_416 ();
 sg13g2_fill_8 FILLER_0_50_424 ();
 sg13g2_fill_8 FILLER_0_50_432 ();
 sg13g2_fill_8 FILLER_0_50_445 ();
 sg13g2_fill_8 FILLER_0_50_453 ();
 sg13g2_fill_8 FILLER_0_50_461 ();
 sg13g2_fill_8 FILLER_0_50_469 ();
 sg13g2_fill_8 FILLER_0_50_477 ();
 sg13g2_fill_4 FILLER_0_50_485 ();
 sg13g2_fill_1 FILLER_0_50_489 ();
 sg13g2_fill_2 FILLER_0_50_498 ();
 sg13g2_fill_2 FILLER_0_50_508 ();
 sg13g2_fill_8 FILLER_0_50_515 ();
 sg13g2_fill_8 FILLER_0_50_523 ();
 sg13g2_fill_8 FILLER_0_50_531 ();
 sg13g2_fill_8 FILLER_0_50_539 ();
 sg13g2_fill_8 FILLER_0_50_547 ();
 sg13g2_fill_8 FILLER_0_50_555 ();
 sg13g2_fill_8 FILLER_0_50_563 ();
 sg13g2_fill_8 FILLER_0_50_571 ();
 sg13g2_fill_8 FILLER_0_50_579 ();
 sg13g2_fill_8 FILLER_0_50_587 ();
 sg13g2_fill_8 FILLER_0_50_595 ();
 sg13g2_fill_8 FILLER_0_50_603 ();
 sg13g2_fill_8 FILLER_0_50_611 ();
 sg13g2_fill_8 FILLER_0_50_619 ();
 sg13g2_fill_8 FILLER_0_50_627 ();
 sg13g2_fill_8 FILLER_0_50_635 ();
 sg13g2_fill_8 FILLER_0_50_643 ();
 sg13g2_fill_8 FILLER_0_50_651 ();
 sg13g2_fill_8 FILLER_0_50_659 ();
 sg13g2_fill_8 FILLER_0_50_667 ();
 sg13g2_fill_1 FILLER_0_50_675 ();
 sg13g2_fill_8 FILLER_0_50_680 ();
 sg13g2_fill_8 FILLER_0_50_688 ();
 sg13g2_fill_1 FILLER_0_50_696 ();
 sg13g2_fill_2 FILLER_0_50_702 ();
 sg13g2_fill_8 FILLER_0_50_709 ();
 sg13g2_fill_8 FILLER_0_50_717 ();
 sg13g2_fill_2 FILLER_0_50_725 ();
 sg13g2_fill_1 FILLER_0_50_727 ();
 sg13g2_fill_8 FILLER_0_50_733 ();
 sg13g2_fill_4 FILLER_0_50_741 ();
 sg13g2_fill_4 FILLER_0_50_749 ();
 sg13g2_fill_2 FILLER_0_50_757 ();
 sg13g2_fill_2 FILLER_0_50_764 ();
 sg13g2_fill_8 FILLER_0_50_787 ();
 sg13g2_fill_2 FILLER_0_50_795 ();
 sg13g2_fill_1 FILLER_0_50_797 ();
 sg13g2_fill_8 FILLER_0_50_803 ();
 sg13g2_fill_8 FILLER_0_50_811 ();
 sg13g2_fill_2 FILLER_0_50_824 ();
 sg13g2_fill_8 FILLER_0_50_831 ();
 sg13g2_fill_8 FILLER_0_50_839 ();
 sg13g2_fill_8 FILLER_0_50_847 ();
 sg13g2_fill_8 FILLER_0_50_855 ();
 sg13g2_fill_4 FILLER_0_50_863 ();
 sg13g2_fill_2 FILLER_0_50_867 ();
 sg13g2_fill_8 FILLER_0_50_874 ();
 sg13g2_fill_8 FILLER_0_50_882 ();
 sg13g2_fill_8 FILLER_0_50_890 ();
 sg13g2_fill_8 FILLER_0_50_898 ();
 sg13g2_fill_8 FILLER_0_50_906 ();
 sg13g2_fill_4 FILLER_0_50_918 ();
 sg13g2_fill_8 FILLER_0_50_932 ();
 sg13g2_fill_4 FILLER_0_50_940 ();
 sg13g2_fill_1 FILLER_0_50_944 ();
 sg13g2_fill_8 FILLER_0_50_950 ();
 sg13g2_fill_1 FILLER_0_50_958 ();
 sg13g2_fill_8 FILLER_0_50_964 ();
 sg13g2_fill_8 FILLER_0_50_972 ();
 sg13g2_fill_2 FILLER_0_50_980 ();
 sg13g2_fill_1 FILLER_0_50_982 ();
 sg13g2_fill_2 FILLER_0_50_1004 ();
 sg13g2_fill_8 FILLER_0_50_1016 ();
 sg13g2_fill_8 FILLER_0_50_1024 ();
 sg13g2_fill_8 FILLER_0_50_1032 ();
 sg13g2_fill_8 FILLER_0_50_1040 ();
 sg13g2_fill_8 FILLER_0_50_1048 ();
 sg13g2_fill_4 FILLER_0_50_1056 ();
 sg13g2_fill_2 FILLER_0_50_1063 ();
 sg13g2_fill_2 FILLER_0_50_1070 ();
 sg13g2_fill_8 FILLER_0_50_1077 ();
 sg13g2_fill_8 FILLER_0_50_1085 ();
 sg13g2_fill_8 FILLER_0_50_1093 ();
 sg13g2_fill_8 FILLER_0_50_1101 ();
 sg13g2_fill_8 FILLER_0_50_1109 ();
 sg13g2_fill_8 FILLER_0_50_1117 ();
 sg13g2_fill_1 FILLER_0_50_1125 ();
 sg13g2_fill_4 FILLER_0_50_1134 ();
 sg13g2_fill_1 FILLER_0_50_1138 ();
 sg13g2_fill_2 FILLER_0_50_1144 ();
 sg13g2_fill_2 FILLER_0_50_1156 ();
 sg13g2_fill_8 FILLER_0_50_1162 ();
 sg13g2_fill_8 FILLER_0_50_1170 ();
 sg13g2_fill_8 FILLER_0_50_1178 ();
 sg13g2_fill_8 FILLER_0_50_1186 ();
 sg13g2_fill_8 FILLER_0_50_1194 ();
 sg13g2_fill_8 FILLER_0_50_1202 ();
 sg13g2_fill_8 FILLER_0_50_1210 ();
 sg13g2_fill_8 FILLER_0_50_1218 ();
 sg13g2_fill_8 FILLER_0_50_1226 ();
 sg13g2_fill_8 FILLER_0_50_1234 ();
 sg13g2_fill_8 FILLER_0_50_1242 ();
 sg13g2_fill_2 FILLER_0_50_1253 ();
 sg13g2_fill_4 FILLER_0_50_1259 ();
 sg13g2_fill_2 FILLER_0_50_1267 ();
 sg13g2_fill_8 FILLER_0_50_1273 ();
 sg13g2_fill_4 FILLER_0_50_1281 ();
 sg13g2_fill_1 FILLER_0_50_1285 ();
 sg13g2_fill_2 FILLER_0_50_1290 ();
 sg13g2_fill_1 FILLER_0_50_1296 ();
 sg13g2_fill_8 FILLER_0_51_0 ();
 sg13g2_fill_8 FILLER_0_51_8 ();
 sg13g2_fill_8 FILLER_0_51_16 ();
 sg13g2_fill_8 FILLER_0_51_24 ();
 sg13g2_fill_8 FILLER_0_51_32 ();
 sg13g2_fill_8 FILLER_0_51_40 ();
 sg13g2_fill_8 FILLER_0_51_48 ();
 sg13g2_fill_8 FILLER_0_51_56 ();
 sg13g2_fill_8 FILLER_0_51_64 ();
 sg13g2_fill_8 FILLER_0_51_72 ();
 sg13g2_fill_8 FILLER_0_51_80 ();
 sg13g2_fill_8 FILLER_0_51_88 ();
 sg13g2_fill_8 FILLER_0_51_96 ();
 sg13g2_fill_8 FILLER_0_51_104 ();
 sg13g2_fill_8 FILLER_0_51_112 ();
 sg13g2_fill_8 FILLER_0_51_120 ();
 sg13g2_fill_8 FILLER_0_51_128 ();
 sg13g2_fill_8 FILLER_0_51_136 ();
 sg13g2_fill_8 FILLER_0_51_144 ();
 sg13g2_fill_8 FILLER_0_51_152 ();
 sg13g2_fill_8 FILLER_0_51_160 ();
 sg13g2_fill_8 FILLER_0_51_168 ();
 sg13g2_fill_8 FILLER_0_51_176 ();
 sg13g2_fill_8 FILLER_0_51_184 ();
 sg13g2_fill_8 FILLER_0_51_192 ();
 sg13g2_fill_8 FILLER_0_51_200 ();
 sg13g2_fill_8 FILLER_0_51_208 ();
 sg13g2_fill_8 FILLER_0_51_216 ();
 sg13g2_fill_1 FILLER_0_51_224 ();
 sg13g2_fill_2 FILLER_0_51_230 ();
 sg13g2_fill_2 FILLER_0_51_258 ();
 sg13g2_fill_2 FILLER_0_51_281 ();
 sg13g2_fill_4 FILLER_0_51_288 ();
 sg13g2_fill_2 FILLER_0_51_292 ();
 sg13g2_fill_1 FILLER_0_51_294 ();
 sg13g2_fill_2 FILLER_0_51_300 ();
 sg13g2_fill_8 FILLER_0_51_309 ();
 sg13g2_fill_8 FILLER_0_51_317 ();
 sg13g2_fill_4 FILLER_0_51_325 ();
 sg13g2_fill_1 FILLER_0_51_329 ();
 sg13g2_fill_2 FILLER_0_51_356 ();
 sg13g2_fill_8 FILLER_0_51_368 ();
 sg13g2_fill_8 FILLER_0_51_380 ();
 sg13g2_fill_8 FILLER_0_51_388 ();
 sg13g2_fill_4 FILLER_0_51_396 ();
 sg13g2_fill_2 FILLER_0_51_400 ();
 sg13g2_fill_2 FILLER_0_51_428 ();
 sg13g2_fill_2 FILLER_0_51_435 ();
 sg13g2_fill_2 FILLER_0_51_441 ();
 sg13g2_fill_8 FILLER_0_51_448 ();
 sg13g2_fill_8 FILLER_0_51_456 ();
 sg13g2_fill_1 FILLER_0_51_464 ();
 sg13g2_fill_8 FILLER_0_51_470 ();
 sg13g2_fill_8 FILLER_0_51_478 ();
 sg13g2_fill_2 FILLER_0_51_486 ();
 sg13g2_fill_2 FILLER_0_51_493 ();
 sg13g2_fill_2 FILLER_0_51_500 ();
 sg13g2_fill_2 FILLER_0_51_509 ();
 sg13g2_fill_8 FILLER_0_51_516 ();
 sg13g2_fill_8 FILLER_0_51_524 ();
 sg13g2_fill_8 FILLER_0_51_532 ();
 sg13g2_fill_8 FILLER_0_51_540 ();
 sg13g2_fill_2 FILLER_0_51_548 ();
 sg13g2_fill_1 FILLER_0_51_550 ();
 sg13g2_fill_8 FILLER_0_51_556 ();
 sg13g2_fill_8 FILLER_0_51_564 ();
 sg13g2_fill_8 FILLER_0_51_572 ();
 sg13g2_fill_8 FILLER_0_51_580 ();
 sg13g2_fill_8 FILLER_0_51_588 ();
 sg13g2_fill_8 FILLER_0_51_596 ();
 sg13g2_fill_8 FILLER_0_51_604 ();
 sg13g2_fill_2 FILLER_0_51_612 ();
 sg13g2_fill_1 FILLER_0_51_614 ();
 sg13g2_fill_8 FILLER_0_51_625 ();
 sg13g2_fill_8 FILLER_0_51_633 ();
 sg13g2_fill_8 FILLER_0_51_641 ();
 sg13g2_fill_4 FILLER_0_51_649 ();
 sg13g2_fill_1 FILLER_0_51_653 ();
 sg13g2_fill_8 FILLER_0_51_659 ();
 sg13g2_fill_4 FILLER_0_51_667 ();
 sg13g2_fill_2 FILLER_0_51_671 ();
 sg13g2_fill_2 FILLER_0_51_678 ();
 sg13g2_fill_4 FILLER_0_51_684 ();
 sg13g2_fill_1 FILLER_0_51_688 ();
 sg13g2_fill_8 FILLER_0_51_694 ();
 sg13g2_fill_4 FILLER_0_51_702 ();
 sg13g2_fill_2 FILLER_0_51_712 ();
 sg13g2_fill_4 FILLER_0_51_720 ();
 sg13g2_fill_2 FILLER_0_51_724 ();
 sg13g2_fill_1 FILLER_0_51_726 ();
 sg13g2_fill_2 FILLER_0_51_731 ();
 sg13g2_fill_2 FILLER_0_51_759 ();
 sg13g2_fill_2 FILLER_0_51_787 ();
 sg13g2_fill_8 FILLER_0_51_794 ();
 sg13g2_fill_4 FILLER_0_51_802 ();
 sg13g2_fill_2 FILLER_0_51_806 ();
 sg13g2_fill_1 FILLER_0_51_808 ();
 sg13g2_fill_8 FILLER_0_51_813 ();
 sg13g2_fill_8 FILLER_0_51_821 ();
 sg13g2_fill_4 FILLER_0_51_829 ();
 sg13g2_fill_2 FILLER_0_51_833 ();
 sg13g2_fill_8 FILLER_0_51_840 ();
 sg13g2_fill_1 FILLER_0_51_848 ();
 sg13g2_fill_8 FILLER_0_51_854 ();
 sg13g2_fill_2 FILLER_0_51_862 ();
 sg13g2_fill_4 FILLER_0_51_869 ();
 sg13g2_fill_1 FILLER_0_51_873 ();
 sg13g2_fill_2 FILLER_0_51_880 ();
 sg13g2_fill_1 FILLER_0_51_882 ();
 sg13g2_fill_8 FILLER_0_51_887 ();
 sg13g2_fill_2 FILLER_0_51_895 ();
 sg13g2_fill_1 FILLER_0_51_897 ();
 sg13g2_fill_4 FILLER_0_51_908 ();
 sg13g2_fill_2 FILLER_0_51_912 ();
 sg13g2_fill_2 FILLER_0_51_919 ();
 sg13g2_fill_1 FILLER_0_51_921 ();
 sg13g2_fill_2 FILLER_0_51_927 ();
 sg13g2_fill_4 FILLER_0_51_934 ();
 sg13g2_fill_1 FILLER_0_51_938 ();
 sg13g2_fill_2 FILLER_0_51_943 ();
 sg13g2_fill_1 FILLER_0_51_945 ();
 sg13g2_fill_2 FILLER_0_51_950 ();
 sg13g2_fill_2 FILLER_0_51_973 ();
 sg13g2_fill_1 FILLER_0_51_975 ();
 sg13g2_fill_8 FILLER_0_51_997 ();
 sg13g2_fill_1 FILLER_0_51_1005 ();
 sg13g2_fill_2 FILLER_0_51_1016 ();
 sg13g2_fill_8 FILLER_0_51_1039 ();
 sg13g2_fill_8 FILLER_0_51_1047 ();
 sg13g2_fill_4 FILLER_0_51_1055 ();
 sg13g2_fill_2 FILLER_0_51_1064 ();
 sg13g2_fill_2 FILLER_0_51_1071 ();
 sg13g2_fill_8 FILLER_0_51_1078 ();
 sg13g2_fill_8 FILLER_0_51_1086 ();
 sg13g2_fill_8 FILLER_0_51_1094 ();
 sg13g2_fill_8 FILLER_0_51_1102 ();
 sg13g2_fill_8 FILLER_0_51_1110 ();
 sg13g2_fill_4 FILLER_0_51_1118 ();
 sg13g2_fill_2 FILLER_0_51_1122 ();
 sg13g2_fill_2 FILLER_0_51_1129 ();
 sg13g2_fill_1 FILLER_0_51_1131 ();
 sg13g2_fill_2 FILLER_0_51_1140 ();
 sg13g2_fill_2 FILLER_0_51_1147 ();
 sg13g2_fill_8 FILLER_0_51_1154 ();
 sg13g2_fill_2 FILLER_0_51_1167 ();
 sg13g2_fill_4 FILLER_0_51_1174 ();
 sg13g2_fill_2 FILLER_0_51_1178 ();
 sg13g2_fill_2 FILLER_0_51_1185 ();
 sg13g2_fill_2 FILLER_0_51_1195 ();
 sg13g2_fill_1 FILLER_0_51_1197 ();
 sg13g2_fill_2 FILLER_0_51_1202 ();
 sg13g2_fill_8 FILLER_0_51_1208 ();
 sg13g2_fill_8 FILLER_0_51_1216 ();
 sg13g2_fill_8 FILLER_0_51_1224 ();
 sg13g2_fill_8 FILLER_0_51_1232 ();
 sg13g2_fill_4 FILLER_0_51_1240 ();
 sg13g2_fill_2 FILLER_0_51_1244 ();
 sg13g2_fill_1 FILLER_0_51_1246 ();
 sg13g2_fill_4 FILLER_0_51_1253 ();
 sg13g2_fill_1 FILLER_0_51_1257 ();
 sg13g2_fill_4 FILLER_0_51_1263 ();
 sg13g2_fill_8 FILLER_0_51_1272 ();
 sg13g2_fill_8 FILLER_0_51_1284 ();
 sg13g2_fill_4 FILLER_0_51_1292 ();
 sg13g2_fill_1 FILLER_0_51_1296 ();
 sg13g2_fill_8 FILLER_0_52_0 ();
 sg13g2_fill_8 FILLER_0_52_8 ();
 sg13g2_fill_8 FILLER_0_52_16 ();
 sg13g2_fill_8 FILLER_0_52_24 ();
 sg13g2_fill_8 FILLER_0_52_32 ();
 sg13g2_fill_8 FILLER_0_52_40 ();
 sg13g2_fill_8 FILLER_0_52_48 ();
 sg13g2_fill_8 FILLER_0_52_56 ();
 sg13g2_fill_8 FILLER_0_52_64 ();
 sg13g2_fill_8 FILLER_0_52_72 ();
 sg13g2_fill_8 FILLER_0_52_80 ();
 sg13g2_fill_8 FILLER_0_52_88 ();
 sg13g2_fill_8 FILLER_0_52_96 ();
 sg13g2_fill_8 FILLER_0_52_104 ();
 sg13g2_fill_8 FILLER_0_52_112 ();
 sg13g2_fill_8 FILLER_0_52_120 ();
 sg13g2_fill_8 FILLER_0_52_128 ();
 sg13g2_fill_8 FILLER_0_52_136 ();
 sg13g2_fill_8 FILLER_0_52_144 ();
 sg13g2_fill_8 FILLER_0_52_152 ();
 sg13g2_fill_8 FILLER_0_52_160 ();
 sg13g2_fill_8 FILLER_0_52_168 ();
 sg13g2_fill_8 FILLER_0_52_176 ();
 sg13g2_fill_8 FILLER_0_52_184 ();
 sg13g2_fill_8 FILLER_0_52_192 ();
 sg13g2_fill_8 FILLER_0_52_200 ();
 sg13g2_fill_8 FILLER_0_52_208 ();
 sg13g2_fill_8 FILLER_0_52_216 ();
 sg13g2_fill_8 FILLER_0_52_224 ();
 sg13g2_fill_8 FILLER_0_52_232 ();
 sg13g2_fill_8 FILLER_0_52_240 ();
 sg13g2_fill_4 FILLER_0_52_248 ();
 sg13g2_fill_1 FILLER_0_52_252 ();
 sg13g2_fill_8 FILLER_0_52_279 ();
 sg13g2_fill_8 FILLER_0_52_287 ();
 sg13g2_fill_2 FILLER_0_52_295 ();
 sg13g2_fill_2 FILLER_0_52_323 ();
 sg13g2_fill_1 FILLER_0_52_325 ();
 sg13g2_fill_2 FILLER_0_52_331 ();
 sg13g2_fill_2 FILLER_0_52_338 ();
 sg13g2_fill_2 FILLER_0_52_344 ();
 sg13g2_fill_2 FILLER_0_52_372 ();
 sg13g2_fill_2 FILLER_0_52_378 ();
 sg13g2_fill_8 FILLER_0_52_384 ();
 sg13g2_fill_8 FILLER_0_52_392 ();
 sg13g2_fill_4 FILLER_0_52_400 ();
 sg13g2_fill_2 FILLER_0_52_409 ();
 sg13g2_fill_2 FILLER_0_52_415 ();
 sg13g2_fill_2 FILLER_0_52_443 ();
 sg13g2_fill_1 FILLER_0_52_445 ();
 sg13g2_fill_4 FILLER_0_52_458 ();
 sg13g2_fill_4 FILLER_0_52_488 ();
 sg13g2_fill_4 FILLER_0_52_497 ();
 sg13g2_fill_4 FILLER_0_52_509 ();
 sg13g2_fill_2 FILLER_0_52_513 ();
 sg13g2_fill_2 FILLER_0_52_520 ();
 sg13g2_fill_8 FILLER_0_52_527 ();
 sg13g2_fill_8 FILLER_0_52_535 ();
 sg13g2_fill_8 FILLER_0_52_543 ();
 sg13g2_fill_2 FILLER_0_52_551 ();
 sg13g2_fill_1 FILLER_0_52_553 ();
 sg13g2_fill_2 FILLER_0_52_580 ();
 sg13g2_fill_8 FILLER_0_52_586 ();
 sg13g2_fill_8 FILLER_0_52_594 ();
 sg13g2_fill_8 FILLER_0_52_602 ();
 sg13g2_fill_8 FILLER_0_52_610 ();
 sg13g2_fill_8 FILLER_0_52_618 ();
 sg13g2_fill_8 FILLER_0_52_626 ();
 sg13g2_fill_8 FILLER_0_52_634 ();
 sg13g2_fill_4 FILLER_0_52_642 ();
 sg13g2_fill_2 FILLER_0_52_646 ();
 sg13g2_fill_2 FILLER_0_52_674 ();
 sg13g2_fill_2 FILLER_0_52_681 ();
 sg13g2_fill_1 FILLER_0_52_683 ();
 sg13g2_fill_2 FILLER_0_52_688 ();
 sg13g2_fill_2 FILLER_0_52_716 ();
 sg13g2_fill_2 FILLER_0_52_722 ();
 sg13g2_fill_2 FILLER_0_52_729 ();
 sg13g2_fill_4 FILLER_0_52_735 ();
 sg13g2_fill_1 FILLER_0_52_739 ();
 sg13g2_fill_2 FILLER_0_52_744 ();
 sg13g2_fill_2 FILLER_0_52_767 ();
 sg13g2_fill_1 FILLER_0_52_769 ();
 sg13g2_fill_4 FILLER_0_52_773 ();
 sg13g2_fill_1 FILLER_0_52_777 ();
 sg13g2_fill_4 FILLER_0_52_783 ();
 sg13g2_fill_2 FILLER_0_52_787 ();
 sg13g2_fill_1 FILLER_0_52_789 ();
 sg13g2_fill_4 FILLER_0_52_802 ();
 sg13g2_fill_2 FILLER_0_52_806 ();
 sg13g2_fill_1 FILLER_0_52_808 ();
 sg13g2_fill_4 FILLER_0_52_814 ();
 sg13g2_fill_1 FILLER_0_52_818 ();
 sg13g2_fill_8 FILLER_0_52_845 ();
 sg13g2_fill_4 FILLER_0_52_853 ();
 sg13g2_fill_2 FILLER_0_52_857 ();
 sg13g2_fill_1 FILLER_0_52_859 ();
 sg13g2_fill_4 FILLER_0_52_886 ();
 sg13g2_fill_1 FILLER_0_52_890 ();
 sg13g2_fill_2 FILLER_0_52_896 ();
 sg13g2_fill_4 FILLER_0_52_903 ();
 sg13g2_fill_2 FILLER_0_52_907 ();
 sg13g2_fill_2 FILLER_0_52_919 ();
 sg13g2_fill_4 FILLER_0_52_925 ();
 sg13g2_fill_1 FILLER_0_52_929 ();
 sg13g2_fill_2 FILLER_0_52_935 ();
 sg13g2_fill_8 FILLER_0_52_941 ();
 sg13g2_fill_8 FILLER_0_52_949 ();
 sg13g2_fill_8 FILLER_0_52_957 ();
 sg13g2_fill_8 FILLER_0_52_965 ();
 sg13g2_fill_4 FILLER_0_52_973 ();
 sg13g2_fill_8 FILLER_0_52_998 ();
 sg13g2_fill_4 FILLER_0_52_1006 ();
 sg13g2_fill_2 FILLER_0_52_1020 ();
 sg13g2_fill_1 FILLER_0_52_1022 ();
 sg13g2_fill_8 FILLER_0_52_1044 ();
 sg13g2_fill_8 FILLER_0_52_1052 ();
 sg13g2_fill_2 FILLER_0_52_1060 ();
 sg13g2_fill_2 FILLER_0_52_1070 ();
 sg13g2_fill_1 FILLER_0_52_1072 ();
 sg13g2_fill_8 FILLER_0_52_1081 ();
 sg13g2_fill_2 FILLER_0_52_1089 ();
 sg13g2_fill_1 FILLER_0_52_1091 ();
 sg13g2_fill_8 FILLER_0_52_1097 ();
 sg13g2_fill_8 FILLER_0_52_1105 ();
 sg13g2_fill_8 FILLER_0_52_1113 ();
 sg13g2_fill_4 FILLER_0_52_1121 ();
 sg13g2_fill_2 FILLER_0_52_1130 ();
 sg13g2_fill_8 FILLER_0_52_1137 ();
 sg13g2_fill_8 FILLER_0_52_1145 ();
 sg13g2_fill_8 FILLER_0_52_1153 ();
 sg13g2_fill_8 FILLER_0_52_1161 ();
 sg13g2_fill_4 FILLER_0_52_1169 ();
 sg13g2_fill_1 FILLER_0_52_1173 ();
 sg13g2_fill_2 FILLER_0_52_1178 ();
 sg13g2_fill_4 FILLER_0_52_1188 ();
 sg13g2_fill_1 FILLER_0_52_1192 ();
 sg13g2_fill_4 FILLER_0_52_1198 ();
 sg13g2_fill_4 FILLER_0_52_1212 ();
 sg13g2_fill_1 FILLER_0_52_1216 ();
 sg13g2_fill_4 FILLER_0_52_1222 ();
 sg13g2_fill_2 FILLER_0_52_1226 ();
 sg13g2_fill_1 FILLER_0_52_1228 ();
 sg13g2_fill_8 FILLER_0_52_1234 ();
 sg13g2_fill_1 FILLER_0_52_1242 ();
 sg13g2_fill_2 FILLER_0_52_1249 ();
 sg13g2_fill_2 FILLER_0_52_1256 ();
 sg13g2_fill_2 FILLER_0_52_1262 ();
 sg13g2_fill_2 FILLER_0_52_1268 ();
 sg13g2_fill_2 FILLER_0_52_1275 ();
 sg13g2_fill_1 FILLER_0_52_1277 ();
 sg13g2_fill_2 FILLER_0_52_1283 ();
 sg13g2_fill_2 FILLER_0_52_1289 ();
 sg13g2_fill_1 FILLER_0_52_1291 ();
 sg13g2_fill_1 FILLER_0_52_1296 ();
 sg13g2_fill_8 FILLER_0_53_0 ();
 sg13g2_fill_8 FILLER_0_53_8 ();
 sg13g2_fill_8 FILLER_0_53_16 ();
 sg13g2_fill_8 FILLER_0_53_24 ();
 sg13g2_fill_8 FILLER_0_53_32 ();
 sg13g2_fill_8 FILLER_0_53_40 ();
 sg13g2_fill_8 FILLER_0_53_48 ();
 sg13g2_fill_8 FILLER_0_53_56 ();
 sg13g2_fill_8 FILLER_0_53_64 ();
 sg13g2_fill_8 FILLER_0_53_72 ();
 sg13g2_fill_8 FILLER_0_53_80 ();
 sg13g2_fill_8 FILLER_0_53_88 ();
 sg13g2_fill_8 FILLER_0_53_96 ();
 sg13g2_fill_8 FILLER_0_53_104 ();
 sg13g2_fill_8 FILLER_0_53_112 ();
 sg13g2_fill_8 FILLER_0_53_120 ();
 sg13g2_fill_8 FILLER_0_53_128 ();
 sg13g2_fill_8 FILLER_0_53_136 ();
 sg13g2_fill_8 FILLER_0_53_144 ();
 sg13g2_fill_8 FILLER_0_53_152 ();
 sg13g2_fill_8 FILLER_0_53_160 ();
 sg13g2_fill_8 FILLER_0_53_168 ();
 sg13g2_fill_8 FILLER_0_53_176 ();
 sg13g2_fill_8 FILLER_0_53_184 ();
 sg13g2_fill_8 FILLER_0_53_192 ();
 sg13g2_fill_8 FILLER_0_53_200 ();
 sg13g2_fill_8 FILLER_0_53_208 ();
 sg13g2_fill_8 FILLER_0_53_216 ();
 sg13g2_fill_8 FILLER_0_53_224 ();
 sg13g2_fill_8 FILLER_0_53_232 ();
 sg13g2_fill_8 FILLER_0_53_240 ();
 sg13g2_fill_1 FILLER_0_53_248 ();
 sg13g2_fill_4 FILLER_0_53_254 ();
 sg13g2_fill_1 FILLER_0_53_258 ();
 sg13g2_fill_8 FILLER_0_53_263 ();
 sg13g2_fill_4 FILLER_0_53_271 ();
 sg13g2_fill_2 FILLER_0_53_280 ();
 sg13g2_fill_8 FILLER_0_53_286 ();
 sg13g2_fill_4 FILLER_0_53_294 ();
 sg13g2_fill_2 FILLER_0_53_298 ();
 sg13g2_fill_8 FILLER_0_53_305 ();
 sg13g2_fill_2 FILLER_0_53_313 ();
 sg13g2_fill_1 FILLER_0_53_315 ();
 sg13g2_fill_2 FILLER_0_53_320 ();
 sg13g2_fill_8 FILLER_0_53_327 ();
 sg13g2_fill_4 FILLER_0_53_335 ();
 sg13g2_fill_1 FILLER_0_53_339 ();
 sg13g2_fill_8 FILLER_0_53_345 ();
 sg13g2_fill_8 FILLER_0_53_353 ();
 sg13g2_fill_8 FILLER_0_53_361 ();
 sg13g2_fill_2 FILLER_0_53_374 ();
 sg13g2_fill_1 FILLER_0_53_376 ();
 sg13g2_fill_2 FILLER_0_53_403 ();
 sg13g2_fill_8 FILLER_0_53_410 ();
 sg13g2_fill_2 FILLER_0_53_418 ();
 sg13g2_fill_1 FILLER_0_53_420 ();
 sg13g2_fill_8 FILLER_0_53_442 ();
 sg13g2_fill_8 FILLER_0_53_450 ();
 sg13g2_fill_2 FILLER_0_53_458 ();
 sg13g2_fill_1 FILLER_0_53_460 ();
 sg13g2_fill_2 FILLER_0_53_466 ();
 sg13g2_fill_8 FILLER_0_53_472 ();
 sg13g2_fill_4 FILLER_0_53_480 ();
 sg13g2_fill_2 FILLER_0_53_484 ();
 sg13g2_fill_4 FILLER_0_53_490 ();
 sg13g2_fill_1 FILLER_0_53_494 ();
 sg13g2_fill_4 FILLER_0_53_521 ();
 sg13g2_fill_2 FILLER_0_53_525 ();
 sg13g2_fill_8 FILLER_0_53_532 ();
 sg13g2_fill_8 FILLER_0_53_540 ();
 sg13g2_fill_2 FILLER_0_53_552 ();
 sg13g2_fill_4 FILLER_0_53_559 ();
 sg13g2_fill_2 FILLER_0_53_567 ();
 sg13g2_fill_1 FILLER_0_53_569 ();
 sg13g2_fill_8 FILLER_0_53_596 ();
 sg13g2_fill_2 FILLER_0_53_604 ();
 sg13g2_fill_1 FILLER_0_53_606 ();
 sg13g2_fill_2 FILLER_0_53_633 ();
 sg13g2_fill_1 FILLER_0_53_635 ();
 sg13g2_fill_4 FILLER_0_53_641 ();
 sg13g2_fill_1 FILLER_0_53_645 ();
 sg13g2_fill_2 FILLER_0_53_652 ();
 sg13g2_fill_8 FILLER_0_53_659 ();
 sg13g2_fill_4 FILLER_0_53_667 ();
 sg13g2_fill_4 FILLER_0_53_677 ();
 sg13g2_fill_2 FILLER_0_53_681 ();
 sg13g2_fill_1 FILLER_0_53_683 ();
 sg13g2_fill_8 FILLER_0_53_688 ();
 sg13g2_fill_8 FILLER_0_53_696 ();
 sg13g2_fill_2 FILLER_0_53_730 ();
 sg13g2_fill_8 FILLER_0_53_737 ();
 sg13g2_fill_2 FILLER_0_53_745 ();
 sg13g2_fill_1 FILLER_0_53_747 ();
 sg13g2_fill_8 FILLER_0_53_753 ();
 sg13g2_fill_4 FILLER_0_53_761 ();
 sg13g2_fill_2 FILLER_0_53_765 ();
 sg13g2_fill_8 FILLER_0_53_773 ();
 sg13g2_fill_8 FILLER_0_53_781 ();
 sg13g2_fill_8 FILLER_0_53_789 ();
 sg13g2_fill_8 FILLER_0_53_797 ();
 sg13g2_fill_4 FILLER_0_53_805 ();
 sg13g2_fill_1 FILLER_0_53_809 ();
 sg13g2_fill_2 FILLER_0_53_815 ();
 sg13g2_fill_1 FILLER_0_53_817 ();
 sg13g2_fill_2 FILLER_0_53_844 ();
 sg13g2_fill_1 FILLER_0_53_846 ();
 sg13g2_fill_2 FILLER_0_53_868 ();
 sg13g2_fill_1 FILLER_0_53_870 ();
 sg13g2_fill_8 FILLER_0_53_879 ();
 sg13g2_fill_8 FILLER_0_53_887 ();
 sg13g2_fill_8 FILLER_0_53_895 ();
 sg13g2_fill_8 FILLER_0_53_903 ();
 sg13g2_fill_2 FILLER_0_53_921 ();
 sg13g2_fill_8 FILLER_0_53_928 ();
 sg13g2_fill_8 FILLER_0_53_936 ();
 sg13g2_fill_2 FILLER_0_53_944 ();
 sg13g2_fill_8 FILLER_0_53_951 ();
 sg13g2_fill_8 FILLER_0_53_959 ();
 sg13g2_fill_8 FILLER_0_53_967 ();
 sg13g2_fill_8 FILLER_0_53_975 ();
 sg13g2_fill_2 FILLER_0_53_983 ();
 sg13g2_fill_2 FILLER_0_53_995 ();
 sg13g2_fill_8 FILLER_0_53_1004 ();
 sg13g2_fill_8 FILLER_0_53_1012 ();
 sg13g2_fill_8 FILLER_0_53_1020 ();
 sg13g2_fill_8 FILLER_0_53_1028 ();
 sg13g2_fill_8 FILLER_0_53_1036 ();
 sg13g2_fill_8 FILLER_0_53_1044 ();
 sg13g2_fill_8 FILLER_0_53_1052 ();
 sg13g2_fill_8 FILLER_0_53_1060 ();
 sg13g2_fill_2 FILLER_0_53_1068 ();
 sg13g2_fill_1 FILLER_0_53_1070 ();
 sg13g2_fill_8 FILLER_0_53_1076 ();
 sg13g2_fill_4 FILLER_0_53_1084 ();
 sg13g2_fill_2 FILLER_0_53_1088 ();
 sg13g2_fill_1 FILLER_0_53_1090 ();
 sg13g2_fill_2 FILLER_0_53_1095 ();
 sg13g2_fill_2 FILLER_0_53_1102 ();
 sg13g2_fill_8 FILLER_0_53_1109 ();
 sg13g2_fill_8 FILLER_0_53_1117 ();
 sg13g2_fill_4 FILLER_0_53_1125 ();
 sg13g2_fill_1 FILLER_0_53_1129 ();
 sg13g2_fill_2 FILLER_0_53_1135 ();
 sg13g2_fill_8 FILLER_0_53_1142 ();
 sg13g2_fill_8 FILLER_0_53_1150 ();
 sg13g2_fill_8 FILLER_0_53_1158 ();
 sg13g2_fill_4 FILLER_0_53_1166 ();
 sg13g2_fill_2 FILLER_0_53_1178 ();
 sg13g2_fill_2 FILLER_0_53_1185 ();
 sg13g2_fill_1 FILLER_0_53_1187 ();
 sg13g2_fill_4 FILLER_0_53_1192 ();
 sg13g2_fill_2 FILLER_0_53_1200 ();
 sg13g2_fill_1 FILLER_0_53_1202 ();
 sg13g2_fill_4 FILLER_0_53_1208 ();
 sg13g2_fill_2 FILLER_0_53_1220 ();
 sg13g2_fill_8 FILLER_0_53_1227 ();
 sg13g2_fill_8 FILLER_0_53_1235 ();
 sg13g2_fill_8 FILLER_0_53_1243 ();
 sg13g2_fill_2 FILLER_0_53_1251 ();
 sg13g2_fill_2 FILLER_0_53_1258 ();
 sg13g2_fill_2 FILLER_0_53_1264 ();
 sg13g2_fill_2 FILLER_0_53_1271 ();
 sg13g2_fill_2 FILLER_0_53_1278 ();
 sg13g2_fill_8 FILLER_0_53_1284 ();
 sg13g2_fill_1 FILLER_0_53_1296 ();
 sg13g2_fill_8 FILLER_0_54_0 ();
 sg13g2_fill_8 FILLER_0_54_8 ();
 sg13g2_fill_8 FILLER_0_54_16 ();
 sg13g2_fill_8 FILLER_0_54_24 ();
 sg13g2_fill_8 FILLER_0_54_32 ();
 sg13g2_fill_8 FILLER_0_54_40 ();
 sg13g2_fill_8 FILLER_0_54_48 ();
 sg13g2_fill_8 FILLER_0_54_56 ();
 sg13g2_fill_8 FILLER_0_54_64 ();
 sg13g2_fill_8 FILLER_0_54_72 ();
 sg13g2_fill_8 FILLER_0_54_80 ();
 sg13g2_fill_8 FILLER_0_54_88 ();
 sg13g2_fill_8 FILLER_0_54_96 ();
 sg13g2_fill_8 FILLER_0_54_104 ();
 sg13g2_fill_8 FILLER_0_54_112 ();
 sg13g2_fill_8 FILLER_0_54_120 ();
 sg13g2_fill_8 FILLER_0_54_128 ();
 sg13g2_fill_8 FILLER_0_54_136 ();
 sg13g2_fill_8 FILLER_0_54_144 ();
 sg13g2_fill_8 FILLER_0_54_152 ();
 sg13g2_fill_8 FILLER_0_54_160 ();
 sg13g2_fill_8 FILLER_0_54_168 ();
 sg13g2_fill_8 FILLER_0_54_176 ();
 sg13g2_fill_8 FILLER_0_54_184 ();
 sg13g2_fill_8 FILLER_0_54_192 ();
 sg13g2_fill_8 FILLER_0_54_200 ();
 sg13g2_fill_8 FILLER_0_54_208 ();
 sg13g2_fill_4 FILLER_0_54_216 ();
 sg13g2_fill_2 FILLER_0_54_220 ();
 sg13g2_fill_1 FILLER_0_54_222 ();
 sg13g2_fill_2 FILLER_0_54_228 ();
 sg13g2_fill_8 FILLER_0_54_234 ();
 sg13g2_fill_8 FILLER_0_54_242 ();
 sg13g2_fill_8 FILLER_0_54_250 ();
 sg13g2_fill_8 FILLER_0_54_258 ();
 sg13g2_fill_8 FILLER_0_54_266 ();
 sg13g2_fill_4 FILLER_0_54_274 ();
 sg13g2_fill_4 FILLER_0_54_304 ();
 sg13g2_fill_1 FILLER_0_54_308 ();
 sg13g2_fill_4 FILLER_0_54_314 ();
 sg13g2_fill_2 FILLER_0_54_318 ();
 sg13g2_fill_8 FILLER_0_54_325 ();
 sg13g2_fill_8 FILLER_0_54_333 ();
 sg13g2_fill_8 FILLER_0_54_341 ();
 sg13g2_fill_8 FILLER_0_54_349 ();
 sg13g2_fill_8 FILLER_0_54_357 ();
 sg13g2_fill_8 FILLER_0_54_365 ();
 sg13g2_fill_8 FILLER_0_54_373 ();
 sg13g2_fill_8 FILLER_0_54_381 ();
 sg13g2_fill_8 FILLER_0_54_389 ();
 sg13g2_fill_2 FILLER_0_54_397 ();
 sg13g2_fill_8 FILLER_0_54_403 ();
 sg13g2_fill_8 FILLER_0_54_411 ();
 sg13g2_fill_8 FILLER_0_54_419 ();
 sg13g2_fill_8 FILLER_0_54_427 ();
 sg13g2_fill_8 FILLER_0_54_445 ();
 sg13g2_fill_8 FILLER_0_54_453 ();
 sg13g2_fill_8 FILLER_0_54_461 ();
 sg13g2_fill_8 FILLER_0_54_469 ();
 sg13g2_fill_4 FILLER_0_54_477 ();
 sg13g2_fill_1 FILLER_0_54_481 ();
 sg13g2_fill_2 FILLER_0_54_487 ();
 sg13g2_fill_8 FILLER_0_54_493 ();
 sg13g2_fill_8 FILLER_0_54_501 ();
 sg13g2_fill_2 FILLER_0_54_509 ();
 sg13g2_fill_1 FILLER_0_54_511 ();
 sg13g2_fill_4 FILLER_0_54_522 ();
 sg13g2_fill_2 FILLER_0_54_526 ();
 sg13g2_fill_2 FILLER_0_54_532 ();
 sg13g2_fill_1 FILLER_0_54_534 ();
 sg13g2_fill_4 FILLER_0_54_540 ();
 sg13g2_fill_1 FILLER_0_54_544 ();
 sg13g2_fill_8 FILLER_0_54_550 ();
 sg13g2_fill_4 FILLER_0_54_558 ();
 sg13g2_fill_2 FILLER_0_54_562 ();
 sg13g2_fill_1 FILLER_0_54_564 ();
 sg13g2_fill_2 FILLER_0_54_570 ();
 sg13g2_fill_2 FILLER_0_54_598 ();
 sg13g2_fill_2 FILLER_0_54_621 ();
 sg13g2_fill_2 FILLER_0_54_628 ();
 sg13g2_fill_8 FILLER_0_54_634 ();
 sg13g2_fill_8 FILLER_0_54_642 ();
 sg13g2_fill_4 FILLER_0_54_650 ();
 sg13g2_fill_2 FILLER_0_54_654 ();
 sg13g2_fill_2 FILLER_0_54_661 ();
 sg13g2_fill_2 FILLER_0_54_667 ();
 sg13g2_fill_1 FILLER_0_54_669 ();
 sg13g2_fill_2 FILLER_0_54_675 ();
 sg13g2_fill_8 FILLER_0_54_683 ();
 sg13g2_fill_8 FILLER_0_54_691 ();
 sg13g2_fill_8 FILLER_0_54_699 ();
 sg13g2_fill_4 FILLER_0_54_707 ();
 sg13g2_fill_2 FILLER_0_54_711 ();
 sg13g2_fill_8 FILLER_0_54_717 ();
 sg13g2_fill_8 FILLER_0_54_725 ();
 sg13g2_fill_8 FILLER_0_54_733 ();
 sg13g2_fill_8 FILLER_0_54_746 ();
 sg13g2_fill_8 FILLER_0_54_754 ();
 sg13g2_fill_8 FILLER_0_54_762 ();
 sg13g2_fill_4 FILLER_0_54_770 ();
 sg13g2_fill_1 FILLER_0_54_774 ();
 sg13g2_fill_8 FILLER_0_54_779 ();
 sg13g2_fill_2 FILLER_0_54_792 ();
 sg13g2_fill_2 FILLER_0_54_799 ();
 sg13g2_fill_8 FILLER_0_54_805 ();
 sg13g2_fill_8 FILLER_0_54_813 ();
 sg13g2_fill_2 FILLER_0_54_821 ();
 sg13g2_fill_2 FILLER_0_54_828 ();
 sg13g2_fill_2 FILLER_0_54_834 ();
 sg13g2_fill_1 FILLER_0_54_836 ();
 sg13g2_fill_8 FILLER_0_54_843 ();
 sg13g2_fill_4 FILLER_0_54_851 ();
 sg13g2_fill_2 FILLER_0_54_855 ();
 sg13g2_fill_2 FILLER_0_54_865 ();
 sg13g2_fill_2 FILLER_0_54_873 ();
 sg13g2_fill_4 FILLER_0_54_880 ();
 sg13g2_fill_2 FILLER_0_54_884 ();
 sg13g2_fill_1 FILLER_0_54_886 ();
 sg13g2_fill_8 FILLER_0_54_892 ();
 sg13g2_fill_4 FILLER_0_54_900 ();
 sg13g2_fill_2 FILLER_0_54_914 ();
 sg13g2_fill_4 FILLER_0_54_920 ();
 sg13g2_fill_1 FILLER_0_54_924 ();
 sg13g2_fill_8 FILLER_0_54_929 ();
 sg13g2_fill_4 FILLER_0_54_937 ();
 sg13g2_fill_2 FILLER_0_54_946 ();
 sg13g2_fill_8 FILLER_0_54_969 ();
 sg13g2_fill_8 FILLER_0_54_981 ();
 sg13g2_fill_2 FILLER_0_54_999 ();
 sg13g2_fill_8 FILLER_0_54_1006 ();
 sg13g2_fill_8 FILLER_0_54_1024 ();
 sg13g2_fill_8 FILLER_0_54_1032 ();
 sg13g2_fill_8 FILLER_0_54_1040 ();
 sg13g2_fill_8 FILLER_0_54_1048 ();
 sg13g2_fill_8 FILLER_0_54_1056 ();
 sg13g2_fill_4 FILLER_0_54_1064 ();
 sg13g2_fill_1 FILLER_0_54_1068 ();
 sg13g2_fill_2 FILLER_0_54_1073 ();
 sg13g2_fill_2 FILLER_0_54_1080 ();
 sg13g2_fill_2 FILLER_0_54_1087 ();
 sg13g2_fill_2 FILLER_0_54_1094 ();
 sg13g2_fill_2 FILLER_0_54_1102 ();
 sg13g2_fill_8 FILLER_0_54_1109 ();
 sg13g2_fill_8 FILLER_0_54_1117 ();
 sg13g2_fill_8 FILLER_0_54_1125 ();
 sg13g2_fill_4 FILLER_0_54_1133 ();
 sg13g2_fill_4 FILLER_0_54_1142 ();
 sg13g2_fill_8 FILLER_0_54_1150 ();
 sg13g2_fill_8 FILLER_0_54_1158 ();
 sg13g2_fill_8 FILLER_0_54_1166 ();
 sg13g2_fill_4 FILLER_0_54_1174 ();
 sg13g2_fill_2 FILLER_0_54_1178 ();
 sg13g2_fill_1 FILLER_0_54_1180 ();
 sg13g2_fill_2 FILLER_0_54_1186 ();
 sg13g2_fill_8 FILLER_0_54_1193 ();
 sg13g2_fill_8 FILLER_0_54_1201 ();
 sg13g2_fill_4 FILLER_0_54_1209 ();
 sg13g2_fill_1 FILLER_0_54_1213 ();
 sg13g2_fill_2 FILLER_0_54_1218 ();
 sg13g2_fill_8 FILLER_0_54_1230 ();
 sg13g2_fill_8 FILLER_0_54_1238 ();
 sg13g2_fill_4 FILLER_0_54_1246 ();
 sg13g2_fill_2 FILLER_0_54_1276 ();
 sg13g2_fill_4 FILLER_0_54_1286 ();
 sg13g2_fill_2 FILLER_0_54_1290 ();
 sg13g2_fill_1 FILLER_0_54_1296 ();
 sg13g2_fill_8 FILLER_0_55_0 ();
 sg13g2_fill_8 FILLER_0_55_8 ();
 sg13g2_fill_8 FILLER_0_55_16 ();
 sg13g2_fill_8 FILLER_0_55_24 ();
 sg13g2_fill_8 FILLER_0_55_32 ();
 sg13g2_fill_8 FILLER_0_55_40 ();
 sg13g2_fill_8 FILLER_0_55_48 ();
 sg13g2_fill_8 FILLER_0_55_56 ();
 sg13g2_fill_8 FILLER_0_55_64 ();
 sg13g2_fill_8 FILLER_0_55_72 ();
 sg13g2_fill_8 FILLER_0_55_80 ();
 sg13g2_fill_8 FILLER_0_55_88 ();
 sg13g2_fill_8 FILLER_0_55_96 ();
 sg13g2_fill_8 FILLER_0_55_104 ();
 sg13g2_fill_8 FILLER_0_55_112 ();
 sg13g2_fill_8 FILLER_0_55_120 ();
 sg13g2_fill_8 FILLER_0_55_128 ();
 sg13g2_fill_8 FILLER_0_55_136 ();
 sg13g2_fill_8 FILLER_0_55_144 ();
 sg13g2_fill_8 FILLER_0_55_152 ();
 sg13g2_fill_8 FILLER_0_55_160 ();
 sg13g2_fill_8 FILLER_0_55_168 ();
 sg13g2_fill_8 FILLER_0_55_176 ();
 sg13g2_fill_8 FILLER_0_55_184 ();
 sg13g2_fill_8 FILLER_0_55_192 ();
 sg13g2_fill_8 FILLER_0_55_200 ();
 sg13g2_fill_2 FILLER_0_55_208 ();
 sg13g2_fill_8 FILLER_0_55_236 ();
 sg13g2_fill_8 FILLER_0_55_244 ();
 sg13g2_fill_8 FILLER_0_55_252 ();
 sg13g2_fill_8 FILLER_0_55_260 ();
 sg13g2_fill_8 FILLER_0_55_268 ();
 sg13g2_fill_8 FILLER_0_55_276 ();
 sg13g2_fill_4 FILLER_0_55_284 ();
 sg13g2_fill_1 FILLER_0_55_288 ();
 sg13g2_fill_2 FILLER_0_55_294 ();
 sg13g2_fill_2 FILLER_0_55_322 ();
 sg13g2_fill_8 FILLER_0_55_328 ();
 sg13g2_fill_8 FILLER_0_55_336 ();
 sg13g2_fill_8 FILLER_0_55_349 ();
 sg13g2_fill_8 FILLER_0_55_357 ();
 sg13g2_fill_8 FILLER_0_55_365 ();
 sg13g2_fill_2 FILLER_0_55_373 ();
 sg13g2_fill_1 FILLER_0_55_375 ();
 sg13g2_fill_4 FILLER_0_55_381 ();
 sg13g2_fill_2 FILLER_0_55_385 ();
 sg13g2_fill_8 FILLER_0_55_391 ();
 sg13g2_fill_8 FILLER_0_55_399 ();
 sg13g2_fill_4 FILLER_0_55_407 ();
 sg13g2_fill_2 FILLER_0_55_411 ();
 sg13g2_fill_1 FILLER_0_55_413 ();
 sg13g2_fill_2 FILLER_0_55_419 ();
 sg13g2_fill_2 FILLER_0_55_427 ();
 sg13g2_fill_8 FILLER_0_55_434 ();
 sg13g2_fill_1 FILLER_0_55_442 ();
 sg13g2_fill_2 FILLER_0_55_448 ();
 sg13g2_fill_8 FILLER_0_55_456 ();
 sg13g2_fill_8 FILLER_0_55_464 ();
 sg13g2_fill_8 FILLER_0_55_472 ();
 sg13g2_fill_1 FILLER_0_55_480 ();
 sg13g2_fill_4 FILLER_0_55_507 ();
 sg13g2_fill_2 FILLER_0_55_511 ();
 sg13g2_fill_1 FILLER_0_55_513 ();
 sg13g2_fill_4 FILLER_0_55_540 ();
 sg13g2_fill_2 FILLER_0_55_544 ();
 sg13g2_fill_8 FILLER_0_55_550 ();
 sg13g2_fill_8 FILLER_0_55_558 ();
 sg13g2_fill_4 FILLER_0_55_566 ();
 sg13g2_fill_2 FILLER_0_55_570 ();
 sg13g2_fill_2 FILLER_0_55_577 ();
 sg13g2_fill_1 FILLER_0_55_579 ();
 sg13g2_fill_2 FILLER_0_55_584 ();
 sg13g2_fill_2 FILLER_0_55_591 ();
 sg13g2_fill_8 FILLER_0_55_614 ();
 sg13g2_fill_1 FILLER_0_55_622 ();
 sg13g2_fill_8 FILLER_0_55_628 ();
 sg13g2_fill_8 FILLER_0_55_636 ();
 sg13g2_fill_8 FILLER_0_55_644 ();
 sg13g2_fill_1 FILLER_0_55_652 ();
 sg13g2_fill_2 FILLER_0_55_679 ();
 sg13g2_fill_2 FILLER_0_55_685 ();
 sg13g2_fill_8 FILLER_0_55_692 ();
 sg13g2_fill_8 FILLER_0_55_700 ();
 sg13g2_fill_8 FILLER_0_55_708 ();
 sg13g2_fill_8 FILLER_0_55_716 ();
 sg13g2_fill_4 FILLER_0_55_724 ();
 sg13g2_fill_2 FILLER_0_55_728 ();
 sg13g2_fill_2 FILLER_0_55_735 ();
 sg13g2_fill_8 FILLER_0_55_741 ();
 sg13g2_fill_4 FILLER_0_55_749 ();
 sg13g2_fill_2 FILLER_0_55_779 ();
 sg13g2_fill_8 FILLER_0_55_802 ();
 sg13g2_fill_8 FILLER_0_55_810 ();
 sg13g2_fill_8 FILLER_0_55_818 ();
 sg13g2_fill_8 FILLER_0_55_826 ();
 sg13g2_fill_8 FILLER_0_55_834 ();
 sg13g2_fill_8 FILLER_0_55_842 ();
 sg13g2_fill_4 FILLER_0_55_850 ();
 sg13g2_fill_2 FILLER_0_55_854 ();
 sg13g2_fill_4 FILLER_0_55_861 ();
 sg13g2_fill_2 FILLER_0_55_865 ();
 sg13g2_fill_8 FILLER_0_55_875 ();
 sg13g2_fill_8 FILLER_0_55_883 ();
 sg13g2_fill_8 FILLER_0_55_891 ();
 sg13g2_fill_8 FILLER_0_55_899 ();
 sg13g2_fill_4 FILLER_0_55_907 ();
 sg13g2_fill_1 FILLER_0_55_911 ();
 sg13g2_fill_2 FILLER_0_55_916 ();
 sg13g2_fill_2 FILLER_0_55_922 ();
 sg13g2_fill_4 FILLER_0_55_928 ();
 sg13g2_fill_2 FILLER_0_55_932 ();
 sg13g2_fill_1 FILLER_0_55_934 ();
 sg13g2_fill_8 FILLER_0_55_945 ();
 sg13g2_fill_8 FILLER_0_55_957 ();
 sg13g2_fill_8 FILLER_0_55_965 ();
 sg13g2_fill_4 FILLER_0_55_973 ();
 sg13g2_fill_2 FILLER_0_55_977 ();
 sg13g2_fill_2 FILLER_0_55_984 ();
 sg13g2_fill_8 FILLER_0_55_1007 ();
 sg13g2_fill_4 FILLER_0_55_1015 ();
 sg13g2_fill_2 FILLER_0_55_1026 ();
 sg13g2_fill_8 FILLER_0_55_1033 ();
 sg13g2_fill_8 FILLER_0_55_1041 ();
 sg13g2_fill_8 FILLER_0_55_1049 ();
 sg13g2_fill_8 FILLER_0_55_1057 ();
 sg13g2_fill_4 FILLER_0_55_1065 ();
 sg13g2_fill_1 FILLER_0_55_1069 ();
 sg13g2_fill_2 FILLER_0_55_1078 ();
 sg13g2_fill_8 FILLER_0_55_1085 ();
 sg13g2_fill_8 FILLER_0_55_1093 ();
 sg13g2_fill_8 FILLER_0_55_1101 ();
 sg13g2_fill_8 FILLER_0_55_1113 ();
 sg13g2_fill_8 FILLER_0_55_1121 ();
 sg13g2_fill_8 FILLER_0_55_1129 ();
 sg13g2_fill_8 FILLER_0_55_1137 ();
 sg13g2_fill_1 FILLER_0_55_1145 ();
 sg13g2_fill_8 FILLER_0_55_1151 ();
 sg13g2_fill_8 FILLER_0_55_1159 ();
 sg13g2_fill_8 FILLER_0_55_1167 ();
 sg13g2_fill_4 FILLER_0_55_1175 ();
 sg13g2_fill_8 FILLER_0_55_1183 ();
 sg13g2_fill_8 FILLER_0_55_1191 ();
 sg13g2_fill_8 FILLER_0_55_1199 ();
 sg13g2_fill_8 FILLER_0_55_1207 ();
 sg13g2_fill_8 FILLER_0_55_1220 ();
 sg13g2_fill_8 FILLER_0_55_1228 ();
 sg13g2_fill_4 FILLER_0_55_1236 ();
 sg13g2_fill_2 FILLER_0_55_1240 ();
 sg13g2_fill_1 FILLER_0_55_1242 ();
 sg13g2_fill_2 FILLER_0_55_1253 ();
 sg13g2_fill_4 FILLER_0_55_1259 ();
 sg13g2_fill_1 FILLER_0_55_1263 ();
 sg13g2_fill_8 FILLER_0_55_1268 ();
 sg13g2_fill_4 FILLER_0_55_1280 ();
 sg13g2_fill_4 FILLER_0_55_1288 ();
 sg13g2_fill_1 FILLER_0_55_1296 ();
 sg13g2_fill_8 FILLER_0_56_0 ();
 sg13g2_fill_8 FILLER_0_56_8 ();
 sg13g2_fill_8 FILLER_0_56_16 ();
 sg13g2_fill_8 FILLER_0_56_24 ();
 sg13g2_fill_8 FILLER_0_56_32 ();
 sg13g2_fill_8 FILLER_0_56_40 ();
 sg13g2_fill_8 FILLER_0_56_48 ();
 sg13g2_fill_8 FILLER_0_56_56 ();
 sg13g2_fill_8 FILLER_0_56_64 ();
 sg13g2_fill_8 FILLER_0_56_72 ();
 sg13g2_fill_8 FILLER_0_56_80 ();
 sg13g2_fill_8 FILLER_0_56_88 ();
 sg13g2_fill_8 FILLER_0_56_96 ();
 sg13g2_fill_8 FILLER_0_56_104 ();
 sg13g2_fill_8 FILLER_0_56_112 ();
 sg13g2_fill_8 FILLER_0_56_120 ();
 sg13g2_fill_8 FILLER_0_56_128 ();
 sg13g2_fill_8 FILLER_0_56_136 ();
 sg13g2_fill_8 FILLER_0_56_144 ();
 sg13g2_fill_8 FILLER_0_56_152 ();
 sg13g2_fill_8 FILLER_0_56_160 ();
 sg13g2_fill_8 FILLER_0_56_168 ();
 sg13g2_fill_8 FILLER_0_56_176 ();
 sg13g2_fill_8 FILLER_0_56_184 ();
 sg13g2_fill_8 FILLER_0_56_192 ();
 sg13g2_fill_8 FILLER_0_56_200 ();
 sg13g2_fill_8 FILLER_0_56_208 ();
 sg13g2_fill_8 FILLER_0_56_216 ();
 sg13g2_fill_8 FILLER_0_56_224 ();
 sg13g2_fill_2 FILLER_0_56_232 ();
 sg13g2_fill_8 FILLER_0_56_255 ();
 sg13g2_fill_4 FILLER_0_56_263 ();
 sg13g2_fill_1 FILLER_0_56_267 ();
 sg13g2_fill_2 FILLER_0_56_273 ();
 sg13g2_fill_8 FILLER_0_56_279 ();
 sg13g2_fill_4 FILLER_0_56_287 ();
 sg13g2_fill_2 FILLER_0_56_291 ();
 sg13g2_fill_2 FILLER_0_56_299 ();
 sg13g2_fill_2 FILLER_0_56_306 ();
 sg13g2_fill_1 FILLER_0_56_308 ();
 sg13g2_fill_2 FILLER_0_56_313 ();
 sg13g2_fill_1 FILLER_0_56_315 ();
 sg13g2_fill_2 FILLER_0_56_326 ();
 sg13g2_fill_2 FILLER_0_56_334 ();
 sg13g2_fill_4 FILLER_0_56_342 ();
 sg13g2_fill_4 FILLER_0_56_352 ();
 sg13g2_fill_2 FILLER_0_56_356 ();
 sg13g2_fill_4 FILLER_0_56_363 ();
 sg13g2_fill_4 FILLER_0_56_393 ();
 sg13g2_fill_2 FILLER_0_56_397 ();
 sg13g2_fill_2 FILLER_0_56_404 ();
 sg13g2_fill_8 FILLER_0_56_432 ();
 sg13g2_fill_2 FILLER_0_56_445 ();
 sg13g2_fill_8 FILLER_0_56_453 ();
 sg13g2_fill_8 FILLER_0_56_461 ();
 sg13g2_fill_1 FILLER_0_56_469 ();
 sg13g2_fill_2 FILLER_0_56_475 ();
 sg13g2_fill_1 FILLER_0_56_477 ();
 sg13g2_fill_4 FILLER_0_56_482 ();
 sg13g2_fill_4 FILLER_0_56_507 ();
 sg13g2_fill_2 FILLER_0_56_511 ();
 sg13g2_fill_1 FILLER_0_56_513 ();
 sg13g2_fill_2 FILLER_0_56_519 ();
 sg13g2_fill_1 FILLER_0_56_521 ();
 sg13g2_fill_4 FILLER_0_56_526 ();
 sg13g2_fill_2 FILLER_0_56_530 ();
 sg13g2_fill_8 FILLER_0_56_553 ();
 sg13g2_fill_8 FILLER_0_56_561 ();
 sg13g2_fill_8 FILLER_0_56_569 ();
 sg13g2_fill_8 FILLER_0_56_577 ();
 sg13g2_fill_8 FILLER_0_56_585 ();
 sg13g2_fill_4 FILLER_0_56_593 ();
 sg13g2_fill_1 FILLER_0_56_597 ();
 sg13g2_fill_8 FILLER_0_56_603 ();
 sg13g2_fill_8 FILLER_0_56_611 ();
 sg13g2_fill_2 FILLER_0_56_619 ();
 sg13g2_fill_1 FILLER_0_56_621 ();
 sg13g2_fill_4 FILLER_0_56_627 ();
 sg13g2_fill_1 FILLER_0_56_631 ();
 sg13g2_fill_8 FILLER_0_56_636 ();
 sg13g2_fill_8 FILLER_0_56_644 ();
 sg13g2_fill_4 FILLER_0_56_652 ();
 sg13g2_fill_2 FILLER_0_56_656 ();
 sg13g2_fill_1 FILLER_0_56_658 ();
 sg13g2_fill_8 FILLER_0_56_664 ();
 sg13g2_fill_2 FILLER_0_56_672 ();
 sg13g2_fill_4 FILLER_0_56_678 ();
 sg13g2_fill_2 FILLER_0_56_687 ();
 sg13g2_fill_1 FILLER_0_56_689 ();
 sg13g2_fill_2 FILLER_0_56_695 ();
 sg13g2_fill_2 FILLER_0_56_702 ();
 sg13g2_fill_2 FILLER_0_56_709 ();
 sg13g2_fill_8 FILLER_0_56_715 ();
 sg13g2_fill_8 FILLER_0_56_723 ();
 sg13g2_fill_8 FILLER_0_56_731 ();
 sg13g2_fill_8 FILLER_0_56_739 ();
 sg13g2_fill_2 FILLER_0_56_747 ();
 sg13g2_fill_2 FILLER_0_56_775 ();
 sg13g2_fill_2 FILLER_0_56_803 ();
 sg13g2_fill_8 FILLER_0_56_831 ();
 sg13g2_fill_8 FILLER_0_56_839 ();
 sg13g2_fill_4 FILLER_0_56_847 ();
 sg13g2_fill_2 FILLER_0_56_851 ();
 sg13g2_fill_1 FILLER_0_56_853 ();
 sg13g2_fill_8 FILLER_0_56_866 ();
 sg13g2_fill_8 FILLER_0_56_874 ();
 sg13g2_fill_8 FILLER_0_56_882 ();
 sg13g2_fill_8 FILLER_0_56_890 ();
 sg13g2_fill_8 FILLER_0_56_898 ();
 sg13g2_fill_8 FILLER_0_56_906 ();
 sg13g2_fill_4 FILLER_0_56_914 ();
 sg13g2_fill_1 FILLER_0_56_918 ();
 sg13g2_fill_2 FILLER_0_56_924 ();
 sg13g2_fill_2 FILLER_0_56_931 ();
 sg13g2_fill_4 FILLER_0_56_937 ();
 sg13g2_fill_1 FILLER_0_56_941 ();
 sg13g2_fill_2 FILLER_0_56_947 ();
 sg13g2_fill_2 FILLER_0_56_953 ();
 sg13g2_fill_1 FILLER_0_56_955 ();
 sg13g2_fill_8 FILLER_0_56_962 ();
 sg13g2_fill_4 FILLER_0_56_975 ();
 sg13g2_fill_2 FILLER_0_56_979 ();
 sg13g2_fill_8 FILLER_0_56_985 ();
 sg13g2_fill_8 FILLER_0_56_993 ();
 sg13g2_fill_1 FILLER_0_56_1001 ();
 sg13g2_fill_8 FILLER_0_56_1007 ();
 sg13g2_fill_4 FILLER_0_56_1015 ();
 sg13g2_fill_2 FILLER_0_56_1019 ();
 sg13g2_fill_8 FILLER_0_56_1025 ();
 sg13g2_fill_8 FILLER_0_56_1041 ();
 sg13g2_fill_8 FILLER_0_56_1049 ();
 sg13g2_fill_8 FILLER_0_56_1057 ();
 sg13g2_fill_2 FILLER_0_56_1065 ();
 sg13g2_fill_1 FILLER_0_56_1067 ();
 sg13g2_fill_2 FILLER_0_56_1072 ();
 sg13g2_fill_8 FILLER_0_56_1079 ();
 sg13g2_fill_8 FILLER_0_56_1087 ();
 sg13g2_fill_8 FILLER_0_56_1095 ();
 sg13g2_fill_4 FILLER_0_56_1103 ();
 sg13g2_fill_2 FILLER_0_56_1111 ();
 sg13g2_fill_4 FILLER_0_56_1119 ();
 sg13g2_fill_8 FILLER_0_56_1128 ();
 sg13g2_fill_2 FILLER_0_56_1141 ();
 sg13g2_fill_8 FILLER_0_56_1151 ();
 sg13g2_fill_2 FILLER_0_56_1159 ();
 sg13g2_fill_8 FILLER_0_56_1165 ();
 sg13g2_fill_8 FILLER_0_56_1173 ();
 sg13g2_fill_4 FILLER_0_56_1181 ();
 sg13g2_fill_1 FILLER_0_56_1185 ();
 sg13g2_fill_2 FILLER_0_56_1192 ();
 sg13g2_fill_8 FILLER_0_56_1199 ();
 sg13g2_fill_8 FILLER_0_56_1207 ();
 sg13g2_fill_8 FILLER_0_56_1215 ();
 sg13g2_fill_2 FILLER_0_56_1223 ();
 sg13g2_fill_1 FILLER_0_56_1225 ();
 sg13g2_fill_8 FILLER_0_56_1234 ();
 sg13g2_fill_4 FILLER_0_56_1242 ();
 sg13g2_fill_2 FILLER_0_56_1251 ();
 sg13g2_fill_8 FILLER_0_56_1258 ();
 sg13g2_fill_1 FILLER_0_56_1266 ();
 sg13g2_fill_4 FILLER_0_56_1271 ();
 sg13g2_fill_1 FILLER_0_56_1275 ();
 sg13g2_fill_2 FILLER_0_56_1280 ();
 sg13g2_fill_2 FILLER_0_56_1286 ();
 sg13g2_fill_4 FILLER_0_56_1292 ();
 sg13g2_fill_1 FILLER_0_56_1296 ();
 sg13g2_fill_8 FILLER_0_57_0 ();
 sg13g2_fill_8 FILLER_0_57_8 ();
 sg13g2_fill_8 FILLER_0_57_16 ();
 sg13g2_fill_8 FILLER_0_57_24 ();
 sg13g2_fill_8 FILLER_0_57_32 ();
 sg13g2_fill_8 FILLER_0_57_40 ();
 sg13g2_fill_8 FILLER_0_57_48 ();
 sg13g2_fill_8 FILLER_0_57_56 ();
 sg13g2_fill_8 FILLER_0_57_64 ();
 sg13g2_fill_8 FILLER_0_57_72 ();
 sg13g2_fill_8 FILLER_0_57_80 ();
 sg13g2_fill_8 FILLER_0_57_88 ();
 sg13g2_fill_8 FILLER_0_57_96 ();
 sg13g2_fill_8 FILLER_0_57_104 ();
 sg13g2_fill_8 FILLER_0_57_112 ();
 sg13g2_fill_8 FILLER_0_57_120 ();
 sg13g2_fill_8 FILLER_0_57_128 ();
 sg13g2_fill_8 FILLER_0_57_136 ();
 sg13g2_fill_8 FILLER_0_57_144 ();
 sg13g2_fill_8 FILLER_0_57_152 ();
 sg13g2_fill_8 FILLER_0_57_160 ();
 sg13g2_fill_8 FILLER_0_57_168 ();
 sg13g2_fill_8 FILLER_0_57_176 ();
 sg13g2_fill_8 FILLER_0_57_184 ();
 sg13g2_fill_8 FILLER_0_57_192 ();
 sg13g2_fill_8 FILLER_0_57_200 ();
 sg13g2_fill_8 FILLER_0_57_208 ();
 sg13g2_fill_8 FILLER_0_57_216 ();
 sg13g2_fill_8 FILLER_0_57_224 ();
 sg13g2_fill_4 FILLER_0_57_258 ();
 sg13g2_fill_2 FILLER_0_57_288 ();
 sg13g2_fill_8 FILLER_0_57_295 ();
 sg13g2_fill_8 FILLER_0_57_303 ();
 sg13g2_fill_8 FILLER_0_57_311 ();
 sg13g2_fill_8 FILLER_0_57_319 ();
 sg13g2_fill_8 FILLER_0_57_327 ();
 sg13g2_fill_1 FILLER_0_57_335 ();
 sg13g2_fill_2 FILLER_0_57_344 ();
 sg13g2_fill_2 FILLER_0_57_372 ();
 sg13g2_fill_8 FILLER_0_57_382 ();
 sg13g2_fill_1 FILLER_0_57_390 ();
 sg13g2_fill_4 FILLER_0_57_401 ();
 sg13g2_fill_2 FILLER_0_57_405 ();
 sg13g2_fill_1 FILLER_0_57_407 ();
 sg13g2_fill_8 FILLER_0_57_412 ();
 sg13g2_fill_8 FILLER_0_57_420 ();
 sg13g2_fill_8 FILLER_0_57_428 ();
 sg13g2_fill_2 FILLER_0_57_436 ();
 sg13g2_fill_1 FILLER_0_57_438 ();
 sg13g2_fill_2 FILLER_0_57_465 ();
 sg13g2_fill_1 FILLER_0_57_467 ();
 sg13g2_fill_8 FILLER_0_57_494 ();
 sg13g2_fill_8 FILLER_0_57_502 ();
 sg13g2_fill_8 FILLER_0_57_510 ();
 sg13g2_fill_8 FILLER_0_57_518 ();
 sg13g2_fill_8 FILLER_0_57_526 ();
 sg13g2_fill_8 FILLER_0_57_534 ();
 sg13g2_fill_8 FILLER_0_57_542 ();
 sg13g2_fill_8 FILLER_0_57_550 ();
 sg13g2_fill_8 FILLER_0_57_558 ();
 sg13g2_fill_8 FILLER_0_57_566 ();
 sg13g2_fill_8 FILLER_0_57_578 ();
 sg13g2_fill_8 FILLER_0_57_586 ();
 sg13g2_fill_8 FILLER_0_57_594 ();
 sg13g2_fill_8 FILLER_0_57_602 ();
 sg13g2_fill_8 FILLER_0_57_610 ();
 sg13g2_fill_2 FILLER_0_57_618 ();
 sg13g2_fill_1 FILLER_0_57_620 ();
 sg13g2_fill_4 FILLER_0_57_647 ();
 sg13g2_fill_2 FILLER_0_57_656 ();
 sg13g2_fill_8 FILLER_0_57_663 ();
 sg13g2_fill_4 FILLER_0_57_676 ();
 sg13g2_fill_2 FILLER_0_57_680 ();
 sg13g2_fill_1 FILLER_0_57_682 ();
 sg13g2_fill_2 FILLER_0_57_688 ();
 sg13g2_fill_2 FILLER_0_57_695 ();
 sg13g2_fill_8 FILLER_0_57_723 ();
 sg13g2_fill_8 FILLER_0_57_736 ();
 sg13g2_fill_1 FILLER_0_57_744 ();
 sg13g2_fill_2 FILLER_0_57_750 ();
 sg13g2_fill_2 FILLER_0_57_756 ();
 sg13g2_fill_1 FILLER_0_57_758 ();
 sg13g2_fill_2 FILLER_0_57_764 ();
 sg13g2_fill_2 FILLER_0_57_770 ();
 sg13g2_fill_2 FILLER_0_57_776 ();
 sg13g2_fill_8 FILLER_0_57_783 ();
 sg13g2_fill_1 FILLER_0_57_791 ();
 sg13g2_fill_2 FILLER_0_57_796 ();
 sg13g2_fill_8 FILLER_0_57_803 ();
 sg13g2_fill_1 FILLER_0_57_811 ();
 sg13g2_fill_8 FILLER_0_57_817 ();
 sg13g2_fill_2 FILLER_0_57_825 ();
 sg13g2_fill_2 FILLER_0_57_831 ();
 sg13g2_fill_2 FILLER_0_57_859 ();
 sg13g2_fill_1 FILLER_0_57_861 ();
 sg13g2_fill_8 FILLER_0_57_868 ();
 sg13g2_fill_2 FILLER_0_57_876 ();
 sg13g2_fill_2 FILLER_0_57_884 ();
 sg13g2_fill_8 FILLER_0_57_890 ();
 sg13g2_fill_8 FILLER_0_57_898 ();
 sg13g2_fill_1 FILLER_0_57_906 ();
 sg13g2_fill_2 FILLER_0_57_917 ();
 sg13g2_fill_8 FILLER_0_57_924 ();
 sg13g2_fill_8 FILLER_0_57_932 ();
 sg13g2_fill_2 FILLER_0_57_940 ();
 sg13g2_fill_2 FILLER_0_57_947 ();
 sg13g2_fill_2 FILLER_0_57_955 ();
 sg13g2_fill_8 FILLER_0_57_963 ();
 sg13g2_fill_4 FILLER_0_57_971 ();
 sg13g2_fill_2 FILLER_0_57_975 ();
 sg13g2_fill_4 FILLER_0_57_987 ();
 sg13g2_fill_2 FILLER_0_57_999 ();
 sg13g2_fill_1 FILLER_0_57_1001 ();
 sg13g2_fill_8 FILLER_0_57_1007 ();
 sg13g2_fill_4 FILLER_0_57_1015 ();
 sg13g2_fill_2 FILLER_0_57_1019 ();
 sg13g2_fill_4 FILLER_0_57_1027 ();
 sg13g2_fill_8 FILLER_0_57_1034 ();
 sg13g2_fill_8 FILLER_0_57_1042 ();
 sg13g2_fill_8 FILLER_0_57_1050 ();
 sg13g2_fill_2 FILLER_0_57_1058 ();
 sg13g2_fill_2 FILLER_0_57_1064 ();
 sg13g2_fill_2 FILLER_0_57_1071 ();
 sg13g2_fill_2 FILLER_0_57_1078 ();
 sg13g2_fill_8 FILLER_0_57_1085 ();
 sg13g2_fill_1 FILLER_0_57_1093 ();
 sg13g2_fill_8 FILLER_0_57_1098 ();
 sg13g2_fill_4 FILLER_0_57_1106 ();
 sg13g2_fill_1 FILLER_0_57_1110 ();
 sg13g2_fill_2 FILLER_0_57_1115 ();
 sg13g2_fill_2 FILLER_0_57_1122 ();
 sg13g2_fill_2 FILLER_0_57_1129 ();
 sg13g2_fill_1 FILLER_0_57_1131 ();
 sg13g2_fill_8 FILLER_0_57_1137 ();
 sg13g2_fill_8 FILLER_0_57_1145 ();
 sg13g2_fill_2 FILLER_0_57_1161 ();
 sg13g2_fill_8 FILLER_0_57_1168 ();
 sg13g2_fill_8 FILLER_0_57_1176 ();
 sg13g2_fill_1 FILLER_0_57_1184 ();
 sg13g2_fill_2 FILLER_0_57_1190 ();
 sg13g2_fill_8 FILLER_0_57_1196 ();
 sg13g2_fill_4 FILLER_0_57_1204 ();
 sg13g2_fill_8 FILLER_0_57_1213 ();
 sg13g2_fill_4 FILLER_0_57_1221 ();
 sg13g2_fill_1 FILLER_0_57_1225 ();
 sg13g2_fill_2 FILLER_0_57_1231 ();
 sg13g2_fill_8 FILLER_0_57_1241 ();
 sg13g2_fill_4 FILLER_0_57_1249 ();
 sg13g2_fill_2 FILLER_0_57_1253 ();
 sg13g2_fill_2 FILLER_0_57_1259 ();
 sg13g2_fill_4 FILLER_0_57_1269 ();
 sg13g2_fill_2 FILLER_0_57_1278 ();
 sg13g2_fill_1 FILLER_0_57_1280 ();
 sg13g2_fill_4 FILLER_0_57_1286 ();
 sg13g2_fill_1 FILLER_0_57_1290 ();
 sg13g2_fill_2 FILLER_0_57_1295 ();
 sg13g2_fill_8 FILLER_0_58_0 ();
 sg13g2_fill_8 FILLER_0_58_8 ();
 sg13g2_fill_8 FILLER_0_58_16 ();
 sg13g2_fill_8 FILLER_0_58_24 ();
 sg13g2_fill_8 FILLER_0_58_32 ();
 sg13g2_fill_8 FILLER_0_58_40 ();
 sg13g2_fill_8 FILLER_0_58_48 ();
 sg13g2_fill_8 FILLER_0_58_56 ();
 sg13g2_fill_8 FILLER_0_58_64 ();
 sg13g2_fill_8 FILLER_0_58_72 ();
 sg13g2_fill_8 FILLER_0_58_80 ();
 sg13g2_fill_8 FILLER_0_58_88 ();
 sg13g2_fill_8 FILLER_0_58_96 ();
 sg13g2_fill_8 FILLER_0_58_104 ();
 sg13g2_fill_8 FILLER_0_58_112 ();
 sg13g2_fill_8 FILLER_0_58_120 ();
 sg13g2_fill_8 FILLER_0_58_128 ();
 sg13g2_fill_8 FILLER_0_58_136 ();
 sg13g2_fill_8 FILLER_0_58_144 ();
 sg13g2_fill_8 FILLER_0_58_152 ();
 sg13g2_fill_8 FILLER_0_58_160 ();
 sg13g2_fill_8 FILLER_0_58_168 ();
 sg13g2_fill_8 FILLER_0_58_176 ();
 sg13g2_fill_8 FILLER_0_58_184 ();
 sg13g2_fill_8 FILLER_0_58_192 ();
 sg13g2_fill_4 FILLER_0_58_200 ();
 sg13g2_fill_2 FILLER_0_58_204 ();
 sg13g2_fill_1 FILLER_0_58_206 ();
 sg13g2_fill_2 FILLER_0_58_233 ();
 sg13g2_fill_1 FILLER_0_58_235 ();
 sg13g2_fill_2 FILLER_0_58_241 ();
 sg13g2_fill_8 FILLER_0_58_247 ();
 sg13g2_fill_8 FILLER_0_58_255 ();
 sg13g2_fill_8 FILLER_0_58_263 ();
 sg13g2_fill_8 FILLER_0_58_271 ();
 sg13g2_fill_8 FILLER_0_58_279 ();
 sg13g2_fill_8 FILLER_0_58_287 ();
 sg13g2_fill_8 FILLER_0_58_295 ();
 sg13g2_fill_8 FILLER_0_58_303 ();
 sg13g2_fill_8 FILLER_0_58_311 ();
 sg13g2_fill_4 FILLER_0_58_319 ();
 sg13g2_fill_2 FILLER_0_58_323 ();
 sg13g2_fill_8 FILLER_0_58_330 ();
 sg13g2_fill_8 FILLER_0_58_338 ();
 sg13g2_fill_8 FILLER_0_58_351 ();
 sg13g2_fill_4 FILLER_0_58_359 ();
 sg13g2_fill_2 FILLER_0_58_363 ();
 sg13g2_fill_1 FILLER_0_58_365 ();
 sg13g2_fill_4 FILLER_0_58_370 ();
 sg13g2_fill_1 FILLER_0_58_374 ();
 sg13g2_fill_8 FILLER_0_58_401 ();
 sg13g2_fill_8 FILLER_0_58_409 ();
 sg13g2_fill_8 FILLER_0_58_417 ();
 sg13g2_fill_8 FILLER_0_58_425 ();
 sg13g2_fill_1 FILLER_0_58_433 ();
 sg13g2_fill_8 FILLER_0_58_439 ();
 sg13g2_fill_8 FILLER_0_58_447 ();
 sg13g2_fill_4 FILLER_0_58_455 ();
 sg13g2_fill_8 FILLER_0_58_463 ();
 sg13g2_fill_2 FILLER_0_58_471 ();
 sg13g2_fill_1 FILLER_0_58_473 ();
 sg13g2_fill_8 FILLER_0_58_479 ();
 sg13g2_fill_4 FILLER_0_58_487 ();
 sg13g2_fill_2 FILLER_0_58_491 ();
 sg13g2_fill_1 FILLER_0_58_493 ();
 sg13g2_fill_8 FILLER_0_58_499 ();
 sg13g2_fill_8 FILLER_0_58_507 ();
 sg13g2_fill_8 FILLER_0_58_515 ();
 sg13g2_fill_8 FILLER_0_58_523 ();
 sg13g2_fill_8 FILLER_0_58_531 ();
 sg13g2_fill_4 FILLER_0_58_539 ();
 sg13g2_fill_1 FILLER_0_58_543 ();
 sg13g2_fill_2 FILLER_0_58_549 ();
 sg13g2_fill_2 FILLER_0_58_577 ();
 sg13g2_fill_8 FILLER_0_58_584 ();
 sg13g2_fill_4 FILLER_0_58_592 ();
 sg13g2_fill_2 FILLER_0_58_596 ();
 sg13g2_fill_1 FILLER_0_58_598 ();
 sg13g2_fill_8 FILLER_0_58_604 ();
 sg13g2_fill_8 FILLER_0_58_612 ();
 sg13g2_fill_8 FILLER_0_58_620 ();
 sg13g2_fill_2 FILLER_0_58_633 ();
 sg13g2_fill_4 FILLER_0_58_639 ();
 sg13g2_fill_1 FILLER_0_58_643 ();
 sg13g2_fill_2 FILLER_0_58_649 ();
 sg13g2_fill_8 FILLER_0_58_656 ();
 sg13g2_fill_2 FILLER_0_58_664 ();
 sg13g2_fill_2 FILLER_0_58_671 ();
 sg13g2_fill_2 FILLER_0_58_699 ();
 sg13g2_fill_1 FILLER_0_58_701 ();
 sg13g2_fill_8 FILLER_0_58_707 ();
 sg13g2_fill_4 FILLER_0_58_715 ();
 sg13g2_fill_1 FILLER_0_58_719 ();
 sg13g2_fill_8 FILLER_0_58_725 ();
 sg13g2_fill_8 FILLER_0_58_733 ();
 sg13g2_fill_8 FILLER_0_58_741 ();
 sg13g2_fill_2 FILLER_0_58_749 ();
 sg13g2_fill_1 FILLER_0_58_751 ();
 sg13g2_fill_8 FILLER_0_58_757 ();
 sg13g2_fill_2 FILLER_0_58_765 ();
 sg13g2_fill_8 FILLER_0_58_777 ();
 sg13g2_fill_2 FILLER_0_58_785 ();
 sg13g2_fill_4 FILLER_0_58_791 ();
 sg13g2_fill_2 FILLER_0_58_795 ();
 sg13g2_fill_4 FILLER_0_58_807 ();
 sg13g2_fill_2 FILLER_0_58_811 ();
 sg13g2_fill_8 FILLER_0_58_817 ();
 sg13g2_fill_4 FILLER_0_58_829 ();
 sg13g2_fill_1 FILLER_0_58_833 ();
 sg13g2_fill_8 FILLER_0_58_839 ();
 sg13g2_fill_8 FILLER_0_58_847 ();
 sg13g2_fill_2 FILLER_0_58_855 ();
 sg13g2_fill_1 FILLER_0_58_857 ();
 sg13g2_fill_4 FILLER_0_58_863 ();
 sg13g2_fill_1 FILLER_0_58_867 ();
 sg13g2_fill_8 FILLER_0_58_894 ();
 sg13g2_fill_8 FILLER_0_58_902 ();
 sg13g2_fill_4 FILLER_0_58_910 ();
 sg13g2_fill_2 FILLER_0_58_918 ();
 sg13g2_fill_2 FILLER_0_58_926 ();
 sg13g2_fill_4 FILLER_0_58_934 ();
 sg13g2_fill_1 FILLER_0_58_938 ();
 sg13g2_fill_8 FILLER_0_58_945 ();
 sg13g2_fill_8 FILLER_0_58_953 ();
 sg13g2_fill_8 FILLER_0_58_961 ();
 sg13g2_fill_8 FILLER_0_58_969 ();
 sg13g2_fill_8 FILLER_0_58_977 ();
 sg13g2_fill_4 FILLER_0_58_989 ();
 sg13g2_fill_2 FILLER_0_58_998 ();
 sg13g2_fill_2 FILLER_0_58_1005 ();
 sg13g2_fill_1 FILLER_0_58_1007 ();
 sg13g2_fill_2 FILLER_0_58_1012 ();
 sg13g2_fill_2 FILLER_0_58_1018 ();
 sg13g2_fill_2 FILLER_0_58_1024 ();
 sg13g2_fill_2 FILLER_0_58_1031 ();
 sg13g2_fill_4 FILLER_0_58_1038 ();
 sg13g2_fill_2 FILLER_0_58_1042 ();
 sg13g2_fill_8 FILLER_0_58_1049 ();
 sg13g2_fill_2 FILLER_0_58_1057 ();
 sg13g2_fill_2 FILLER_0_58_1064 ();
 sg13g2_fill_2 FILLER_0_58_1071 ();
 sg13g2_fill_4 FILLER_0_58_1077 ();
 sg13g2_fill_2 FILLER_0_58_1081 ();
 sg13g2_fill_1 FILLER_0_58_1083 ();
 sg13g2_fill_2 FILLER_0_58_1089 ();
 sg13g2_fill_2 FILLER_0_58_1099 ();
 sg13g2_fill_8 FILLER_0_58_1106 ();
 sg13g2_fill_2 FILLER_0_58_1114 ();
 sg13g2_fill_2 FILLER_0_58_1126 ();
 sg13g2_fill_2 FILLER_0_58_1132 ();
 sg13g2_fill_1 FILLER_0_58_1134 ();
 sg13g2_fill_2 FILLER_0_58_1139 ();
 sg13g2_fill_8 FILLER_0_58_1146 ();
 sg13g2_fill_1 FILLER_0_58_1154 ();
 sg13g2_fill_4 FILLER_0_58_1160 ();
 sg13g2_fill_2 FILLER_0_58_1164 ();
 sg13g2_fill_4 FILLER_0_58_1171 ();
 sg13g2_fill_4 FILLER_0_58_1180 ();
 sg13g2_fill_1 FILLER_0_58_1184 ();
 sg13g2_fill_2 FILLER_0_58_1191 ();
 sg13g2_fill_4 FILLER_0_58_1198 ();
 sg13g2_fill_2 FILLER_0_58_1208 ();
 sg13g2_fill_1 FILLER_0_58_1210 ();
 sg13g2_fill_4 FILLER_0_58_1216 ();
 sg13g2_fill_8 FILLER_0_58_1225 ();
 sg13g2_fill_1 FILLER_0_58_1233 ();
 sg13g2_fill_2 FILLER_0_58_1239 ();
 sg13g2_fill_2 FILLER_0_58_1246 ();
 sg13g2_fill_8 FILLER_0_58_1252 ();
 sg13g2_fill_4 FILLER_0_58_1260 ();
 sg13g2_fill_1 FILLER_0_58_1264 ();
 sg13g2_fill_2 FILLER_0_58_1270 ();
 sg13g2_fill_4 FILLER_0_58_1276 ();
 sg13g2_fill_2 FILLER_0_58_1280 ();
 sg13g2_fill_8 FILLER_0_58_1287 ();
 sg13g2_fill_2 FILLER_0_58_1295 ();
 sg13g2_fill_8 FILLER_0_59_0 ();
 sg13g2_fill_8 FILLER_0_59_8 ();
 sg13g2_fill_8 FILLER_0_59_16 ();
 sg13g2_fill_8 FILLER_0_59_24 ();
 sg13g2_fill_8 FILLER_0_59_32 ();
 sg13g2_fill_8 FILLER_0_59_40 ();
 sg13g2_fill_8 FILLER_0_59_48 ();
 sg13g2_fill_8 FILLER_0_59_56 ();
 sg13g2_fill_8 FILLER_0_59_64 ();
 sg13g2_fill_8 FILLER_0_59_72 ();
 sg13g2_fill_8 FILLER_0_59_80 ();
 sg13g2_fill_8 FILLER_0_59_88 ();
 sg13g2_fill_8 FILLER_0_59_96 ();
 sg13g2_fill_8 FILLER_0_59_104 ();
 sg13g2_fill_8 FILLER_0_59_112 ();
 sg13g2_fill_8 FILLER_0_59_120 ();
 sg13g2_fill_8 FILLER_0_59_128 ();
 sg13g2_fill_8 FILLER_0_59_136 ();
 sg13g2_fill_8 FILLER_0_59_144 ();
 sg13g2_fill_8 FILLER_0_59_152 ();
 sg13g2_fill_8 FILLER_0_59_160 ();
 sg13g2_fill_8 FILLER_0_59_168 ();
 sg13g2_fill_8 FILLER_0_59_176 ();
 sg13g2_fill_8 FILLER_0_59_184 ();
 sg13g2_fill_8 FILLER_0_59_192 ();
 sg13g2_fill_8 FILLER_0_59_200 ();
 sg13g2_fill_4 FILLER_0_59_208 ();
 sg13g2_fill_2 FILLER_0_59_238 ();
 sg13g2_fill_8 FILLER_0_59_261 ();
 sg13g2_fill_4 FILLER_0_59_269 ();
 sg13g2_fill_8 FILLER_0_59_277 ();
 sg13g2_fill_8 FILLER_0_59_285 ();
 sg13g2_fill_8 FILLER_0_59_293 ();
 sg13g2_fill_2 FILLER_0_59_306 ();
 sg13g2_fill_2 FILLER_0_59_313 ();
 sg13g2_fill_8 FILLER_0_59_319 ();
 sg13g2_fill_8 FILLER_0_59_327 ();
 sg13g2_fill_8 FILLER_0_59_335 ();
 sg13g2_fill_8 FILLER_0_59_343 ();
 sg13g2_fill_8 FILLER_0_59_351 ();
 sg13g2_fill_4 FILLER_0_59_359 ();
 sg13g2_fill_4 FILLER_0_59_368 ();
 sg13g2_fill_4 FILLER_0_59_377 ();
 sg13g2_fill_4 FILLER_0_59_385 ();
 sg13g2_fill_8 FILLER_0_59_410 ();
 sg13g2_fill_2 FILLER_0_59_418 ();
 sg13g2_fill_2 FILLER_0_59_424 ();
 sg13g2_fill_8 FILLER_0_59_434 ();
 sg13g2_fill_2 FILLER_0_59_446 ();
 sg13g2_fill_8 FILLER_0_59_453 ();
 sg13g2_fill_8 FILLER_0_59_461 ();
 sg13g2_fill_8 FILLER_0_59_469 ();
 sg13g2_fill_8 FILLER_0_59_477 ();
 sg13g2_fill_8 FILLER_0_59_485 ();
 sg13g2_fill_4 FILLER_0_59_493 ();
 sg13g2_fill_1 FILLER_0_59_497 ();
 sg13g2_fill_2 FILLER_0_59_504 ();
 sg13g2_fill_4 FILLER_0_59_511 ();
 sg13g2_fill_2 FILLER_0_59_515 ();
 sg13g2_fill_1 FILLER_0_59_517 ();
 sg13g2_fill_2 FILLER_0_59_523 ();
 sg13g2_fill_1 FILLER_0_59_525 ();
 sg13g2_fill_8 FILLER_0_59_530 ();
 sg13g2_fill_8 FILLER_0_59_538 ();
 sg13g2_fill_8 FILLER_0_59_546 ();
 sg13g2_fill_4 FILLER_0_59_554 ();
 sg13g2_fill_2 FILLER_0_59_558 ();
 sg13g2_fill_1 FILLER_0_59_560 ();
 sg13g2_fill_2 FILLER_0_59_565 ();
 sg13g2_fill_1 FILLER_0_59_567 ();
 sg13g2_fill_2 FILLER_0_59_594 ();
 sg13g2_fill_2 FILLER_0_59_599 ();
 sg13g2_fill_2 FILLER_0_59_606 ();
 sg13g2_fill_4 FILLER_0_59_613 ();
 sg13g2_fill_1 FILLER_0_59_617 ();
 sg13g2_fill_2 FILLER_0_59_644 ();
 sg13g2_fill_2 FILLER_0_59_650 ();
 sg13g2_fill_4 FILLER_0_59_658 ();
 sg13g2_fill_2 FILLER_0_59_662 ();
 sg13g2_fill_2 FILLER_0_59_672 ();
 sg13g2_fill_8 FILLER_0_59_679 ();
 sg13g2_fill_2 FILLER_0_59_687 ();
 sg13g2_fill_4 FILLER_0_59_695 ();
 sg13g2_fill_2 FILLER_0_59_699 ();
 sg13g2_fill_1 FILLER_0_59_701 ();
 sg13g2_fill_8 FILLER_0_59_707 ();
 sg13g2_fill_8 FILLER_0_59_715 ();
 sg13g2_fill_8 FILLER_0_59_723 ();
 sg13g2_fill_2 FILLER_0_59_736 ();
 sg13g2_fill_2 FILLER_0_59_742 ();
 sg13g2_fill_2 FILLER_0_59_749 ();
 sg13g2_fill_1 FILLER_0_59_751 ();
 sg13g2_fill_8 FILLER_0_59_756 ();
 sg13g2_fill_2 FILLER_0_59_764 ();
 sg13g2_fill_8 FILLER_0_59_771 ();
 sg13g2_fill_4 FILLER_0_59_784 ();
 sg13g2_fill_2 FILLER_0_59_793 ();
 sg13g2_fill_8 FILLER_0_59_799 ();
 sg13g2_fill_8 FILLER_0_59_807 ();
 sg13g2_fill_4 FILLER_0_59_815 ();
 sg13g2_fill_1 FILLER_0_59_819 ();
 sg13g2_fill_2 FILLER_0_59_825 ();
 sg13g2_fill_2 FILLER_0_59_853 ();
 sg13g2_fill_2 FILLER_0_59_860 ();
 sg13g2_fill_2 FILLER_0_59_867 ();
 sg13g2_fill_2 FILLER_0_59_879 ();
 sg13g2_fill_8 FILLER_0_59_886 ();
 sg13g2_fill_8 FILLER_0_59_894 ();
 sg13g2_fill_8 FILLER_0_59_902 ();
 sg13g2_fill_4 FILLER_0_59_910 ();
 sg13g2_fill_1 FILLER_0_59_914 ();
 sg13g2_fill_2 FILLER_0_59_919 ();
 sg13g2_fill_2 FILLER_0_59_927 ();
 sg13g2_fill_1 FILLER_0_59_929 ();
 sg13g2_fill_8 FILLER_0_59_940 ();
 sg13g2_fill_8 FILLER_0_59_948 ();
 sg13g2_fill_8 FILLER_0_59_956 ();
 sg13g2_fill_8 FILLER_0_59_964 ();
 sg13g2_fill_1 FILLER_0_59_972 ();
 sg13g2_fill_4 FILLER_0_59_977 ();
 sg13g2_fill_2 FILLER_0_59_981 ();
 sg13g2_fill_8 FILLER_0_59_987 ();
 sg13g2_fill_2 FILLER_0_59_999 ();
 sg13g2_fill_1 FILLER_0_59_1001 ();
 sg13g2_fill_8 FILLER_0_59_1007 ();
 sg13g2_fill_4 FILLER_0_59_1015 ();
 sg13g2_fill_2 FILLER_0_59_1019 ();
 sg13g2_fill_1 FILLER_0_59_1021 ();
 sg13g2_fill_2 FILLER_0_59_1026 ();
 sg13g2_fill_1 FILLER_0_59_1028 ();
 sg13g2_fill_2 FILLER_0_59_1036 ();
 sg13g2_fill_8 FILLER_0_59_1043 ();
 sg13g2_fill_8 FILLER_0_59_1051 ();
 sg13g2_fill_8 FILLER_0_59_1059 ();
 sg13g2_fill_8 FILLER_0_59_1067 ();
 sg13g2_fill_2 FILLER_0_59_1075 ();
 sg13g2_fill_8 FILLER_0_59_1082 ();
 sg13g2_fill_1 FILLER_0_59_1090 ();
 sg13g2_fill_8 FILLER_0_59_1096 ();
 sg13g2_fill_8 FILLER_0_59_1104 ();
 sg13g2_fill_8 FILLER_0_59_1112 ();
 sg13g2_fill_2 FILLER_0_59_1120 ();
 sg13g2_fill_1 FILLER_0_59_1122 ();
 sg13g2_fill_2 FILLER_0_59_1128 ();
 sg13g2_fill_8 FILLER_0_59_1134 ();
 sg13g2_fill_8 FILLER_0_59_1142 ();
 sg13g2_fill_2 FILLER_0_59_1150 ();
 sg13g2_fill_4 FILLER_0_59_1160 ();
 sg13g2_fill_2 FILLER_0_59_1164 ();
 sg13g2_fill_1 FILLER_0_59_1166 ();
 sg13g2_fill_2 FILLER_0_59_1172 ();
 sg13g2_fill_1 FILLER_0_59_1174 ();
 sg13g2_fill_2 FILLER_0_59_1181 ();
 sg13g2_fill_2 FILLER_0_59_1188 ();
 sg13g2_fill_2 FILLER_0_59_1195 ();
 sg13g2_fill_2 FILLER_0_59_1202 ();
 sg13g2_fill_8 FILLER_0_59_1208 ();
 sg13g2_fill_4 FILLER_0_59_1216 ();
 sg13g2_fill_2 FILLER_0_59_1220 ();
 sg13g2_fill_4 FILLER_0_59_1228 ();
 sg13g2_fill_2 FILLER_0_59_1232 ();
 sg13g2_fill_4 FILLER_0_59_1240 ();
 sg13g2_fill_2 FILLER_0_59_1244 ();
 sg13g2_fill_1 FILLER_0_59_1246 ();
 sg13g2_fill_2 FILLER_0_59_1273 ();
 sg13g2_fill_2 FILLER_0_59_1280 ();
 sg13g2_fill_1 FILLER_0_59_1282 ();
 sg13g2_fill_4 FILLER_0_59_1288 ();
 sg13g2_fill_1 FILLER_0_59_1296 ();
 sg13g2_fill_8 FILLER_0_60_0 ();
 sg13g2_fill_8 FILLER_0_60_8 ();
 sg13g2_fill_8 FILLER_0_60_16 ();
 sg13g2_fill_8 FILLER_0_60_24 ();
 sg13g2_fill_8 FILLER_0_60_32 ();
 sg13g2_fill_8 FILLER_0_60_40 ();
 sg13g2_fill_8 FILLER_0_60_48 ();
 sg13g2_fill_8 FILLER_0_60_56 ();
 sg13g2_fill_8 FILLER_0_60_64 ();
 sg13g2_fill_8 FILLER_0_60_72 ();
 sg13g2_fill_8 FILLER_0_60_80 ();
 sg13g2_fill_8 FILLER_0_60_88 ();
 sg13g2_fill_8 FILLER_0_60_96 ();
 sg13g2_fill_8 FILLER_0_60_104 ();
 sg13g2_fill_8 FILLER_0_60_112 ();
 sg13g2_fill_8 FILLER_0_60_120 ();
 sg13g2_fill_8 FILLER_0_60_128 ();
 sg13g2_fill_8 FILLER_0_60_136 ();
 sg13g2_fill_8 FILLER_0_60_144 ();
 sg13g2_fill_8 FILLER_0_60_152 ();
 sg13g2_fill_8 FILLER_0_60_160 ();
 sg13g2_fill_8 FILLER_0_60_168 ();
 sg13g2_fill_8 FILLER_0_60_176 ();
 sg13g2_fill_8 FILLER_0_60_184 ();
 sg13g2_fill_8 FILLER_0_60_192 ();
 sg13g2_fill_8 FILLER_0_60_200 ();
 sg13g2_fill_4 FILLER_0_60_208 ();
 sg13g2_fill_2 FILLER_0_60_212 ();
 sg13g2_fill_1 FILLER_0_60_214 ();
 sg13g2_fill_2 FILLER_0_60_220 ();
 sg13g2_fill_2 FILLER_0_60_226 ();
 sg13g2_fill_8 FILLER_0_60_232 ();
 sg13g2_fill_8 FILLER_0_60_240 ();
 sg13g2_fill_8 FILLER_0_60_248 ();
 sg13g2_fill_4 FILLER_0_60_256 ();
 sg13g2_fill_4 FILLER_0_60_267 ();
 sg13g2_fill_4 FILLER_0_60_277 ();
 sg13g2_fill_2 FILLER_0_60_287 ();
 sg13g2_fill_2 FILLER_0_60_294 ();
 sg13g2_fill_2 FILLER_0_60_322 ();
 sg13g2_fill_8 FILLER_0_60_345 ();
 sg13g2_fill_2 FILLER_0_60_353 ();
 sg13g2_fill_8 FILLER_0_60_360 ();
 sg13g2_fill_8 FILLER_0_60_368 ();
 sg13g2_fill_1 FILLER_0_60_376 ();
 sg13g2_fill_8 FILLER_0_60_381 ();
 sg13g2_fill_8 FILLER_0_60_389 ();
 sg13g2_fill_8 FILLER_0_60_397 ();
 sg13g2_fill_2 FILLER_0_60_405 ();
 sg13g2_fill_1 FILLER_0_60_407 ();
 sg13g2_fill_8 FILLER_0_60_412 ();
 sg13g2_fill_4 FILLER_0_60_420 ();
 sg13g2_fill_2 FILLER_0_60_424 ();
 sg13g2_fill_4 FILLER_0_60_430 ();
 sg13g2_fill_2 FILLER_0_60_439 ();
 sg13g2_fill_8 FILLER_0_60_467 ();
 sg13g2_fill_4 FILLER_0_60_475 ();
 sg13g2_fill_2 FILLER_0_60_479 ();
 sg13g2_fill_4 FILLER_0_60_486 ();
 sg13g2_fill_1 FILLER_0_60_490 ();
 sg13g2_fill_8 FILLER_0_60_495 ();
 sg13g2_fill_1 FILLER_0_60_503 ();
 sg13g2_fill_8 FILLER_0_60_510 ();
 sg13g2_fill_8 FILLER_0_60_544 ();
 sg13g2_fill_8 FILLER_0_60_552 ();
 sg13g2_fill_2 FILLER_0_60_560 ();
 sg13g2_fill_2 FILLER_0_60_567 ();
 sg13g2_fill_2 FILLER_0_60_574 ();
 sg13g2_fill_2 FILLER_0_60_586 ();
 sg13g2_fill_4 FILLER_0_60_593 ();
 sg13g2_fill_2 FILLER_0_60_597 ();
 sg13g2_fill_2 FILLER_0_60_605 ();
 sg13g2_fill_8 FILLER_0_60_613 ();
 sg13g2_fill_8 FILLER_0_60_621 ();
 sg13g2_fill_8 FILLER_0_60_629 ();
 sg13g2_fill_1 FILLER_0_60_637 ();
 sg13g2_fill_2 FILLER_0_60_648 ();
 sg13g2_fill_4 FILLER_0_60_655 ();
 sg13g2_fill_2 FILLER_0_60_667 ();
 sg13g2_fill_1 FILLER_0_60_669 ();
 sg13g2_fill_8 FILLER_0_60_675 ();
 sg13g2_fill_4 FILLER_0_60_683 ();
 sg13g2_fill_2 FILLER_0_60_687 ();
 sg13g2_fill_1 FILLER_0_60_689 ();
 sg13g2_fill_8 FILLER_0_60_694 ();
 sg13g2_fill_1 FILLER_0_60_702 ();
 sg13g2_fill_8 FILLER_0_60_711 ();
 sg13g2_fill_8 FILLER_0_60_719 ();
 sg13g2_fill_1 FILLER_0_60_727 ();
 sg13g2_fill_2 FILLER_0_60_754 ();
 sg13g2_fill_2 FILLER_0_60_766 ();
 sg13g2_fill_2 FILLER_0_60_773 ();
 sg13g2_fill_4 FILLER_0_60_779 ();
 sg13g2_fill_4 FILLER_0_60_789 ();
 sg13g2_fill_2 FILLER_0_60_793 ();
 sg13g2_fill_1 FILLER_0_60_795 ();
 sg13g2_fill_4 FILLER_0_60_801 ();
 sg13g2_fill_8 FILLER_0_60_809 ();
 sg13g2_fill_8 FILLER_0_60_817 ();
 sg13g2_fill_4 FILLER_0_60_825 ();
 sg13g2_fill_2 FILLER_0_60_829 ();
 sg13g2_fill_1 FILLER_0_60_831 ();
 sg13g2_fill_8 FILLER_0_60_837 ();
 sg13g2_fill_8 FILLER_0_60_845 ();
 sg13g2_fill_8 FILLER_0_60_853 ();
 sg13g2_fill_8 FILLER_0_60_861 ();
 sg13g2_fill_8 FILLER_0_60_869 ();
 sg13g2_fill_8 FILLER_0_60_877 ();
 sg13g2_fill_8 FILLER_0_60_885 ();
 sg13g2_fill_2 FILLER_0_60_893 ();
 sg13g2_fill_1 FILLER_0_60_895 ();
 sg13g2_fill_2 FILLER_0_60_900 ();
 sg13g2_fill_2 FILLER_0_60_907 ();
 sg13g2_fill_8 FILLER_0_60_914 ();
 sg13g2_fill_4 FILLER_0_60_922 ();
 sg13g2_fill_2 FILLER_0_60_926 ();
 sg13g2_fill_8 FILLER_0_60_938 ();
 sg13g2_fill_2 FILLER_0_60_946 ();
 sg13g2_fill_8 FILLER_0_60_952 ();
 sg13g2_fill_8 FILLER_0_60_960 ();
 sg13g2_fill_1 FILLER_0_60_968 ();
 sg13g2_fill_8 FILLER_0_60_974 ();
 sg13g2_fill_2 FILLER_0_60_987 ();
 sg13g2_fill_2 FILLER_0_60_995 ();
 sg13g2_fill_4 FILLER_0_60_1002 ();
 sg13g2_fill_2 FILLER_0_60_1006 ();
 sg13g2_fill_2 FILLER_0_60_1013 ();
 sg13g2_fill_4 FILLER_0_60_1020 ();
 sg13g2_fill_1 FILLER_0_60_1024 ();
 sg13g2_fill_4 FILLER_0_60_1031 ();
 sg13g2_fill_2 FILLER_0_60_1035 ();
 sg13g2_fill_1 FILLER_0_60_1037 ();
 sg13g2_fill_2 FILLER_0_60_1045 ();
 sg13g2_fill_8 FILLER_0_60_1051 ();
 sg13g2_fill_8 FILLER_0_60_1059 ();
 sg13g2_fill_4 FILLER_0_60_1067 ();
 sg13g2_fill_1 FILLER_0_60_1071 ();
 sg13g2_fill_2 FILLER_0_60_1077 ();
 sg13g2_fill_8 FILLER_0_60_1089 ();
 sg13g2_fill_8 FILLER_0_60_1097 ();
 sg13g2_fill_4 FILLER_0_60_1105 ();
 sg13g2_fill_2 FILLER_0_60_1116 ();
 sg13g2_fill_4 FILLER_0_60_1123 ();
 sg13g2_fill_1 FILLER_0_60_1127 ();
 sg13g2_fill_2 FILLER_0_60_1132 ();
 sg13g2_fill_8 FILLER_0_60_1139 ();
 sg13g2_fill_8 FILLER_0_60_1147 ();
 sg13g2_fill_4 FILLER_0_60_1155 ();
 sg13g2_fill_1 FILLER_0_60_1159 ();
 sg13g2_fill_2 FILLER_0_60_1165 ();
 sg13g2_fill_1 FILLER_0_60_1167 ();
 sg13g2_fill_2 FILLER_0_60_1176 ();
 sg13g2_fill_1 FILLER_0_60_1178 ();
 sg13g2_fill_8 FILLER_0_60_1184 ();
 sg13g2_fill_8 FILLER_0_60_1192 ();
 sg13g2_fill_8 FILLER_0_60_1200 ();
 sg13g2_fill_8 FILLER_0_60_1208 ();
 sg13g2_fill_2 FILLER_0_60_1216 ();
 sg13g2_fill_1 FILLER_0_60_1218 ();
 sg13g2_fill_2 FILLER_0_60_1223 ();
 sg13g2_fill_4 FILLER_0_60_1230 ();
 sg13g2_fill_2 FILLER_0_60_1234 ();
 sg13g2_fill_8 FILLER_0_60_1241 ();
 sg13g2_fill_8 FILLER_0_60_1253 ();
 sg13g2_fill_8 FILLER_0_60_1265 ();
 sg13g2_fill_4 FILLER_0_60_1273 ();
 sg13g2_fill_2 FILLER_0_60_1277 ();
 sg13g2_fill_4 FILLER_0_60_1283 ();
 sg13g2_fill_1 FILLER_0_60_1287 ();
 sg13g2_fill_4 FILLER_0_60_1292 ();
 sg13g2_fill_1 FILLER_0_60_1296 ();
 sg13g2_fill_8 FILLER_0_61_0 ();
 sg13g2_fill_8 FILLER_0_61_8 ();
 sg13g2_fill_8 FILLER_0_61_16 ();
 sg13g2_fill_8 FILLER_0_61_24 ();
 sg13g2_fill_8 FILLER_0_61_32 ();
 sg13g2_fill_8 FILLER_0_61_40 ();
 sg13g2_fill_8 FILLER_0_61_48 ();
 sg13g2_fill_8 FILLER_0_61_56 ();
 sg13g2_fill_8 FILLER_0_61_64 ();
 sg13g2_fill_8 FILLER_0_61_72 ();
 sg13g2_fill_8 FILLER_0_61_80 ();
 sg13g2_fill_8 FILLER_0_61_88 ();
 sg13g2_fill_8 FILLER_0_61_96 ();
 sg13g2_fill_8 FILLER_0_61_104 ();
 sg13g2_fill_8 FILLER_0_61_112 ();
 sg13g2_fill_8 FILLER_0_61_120 ();
 sg13g2_fill_8 FILLER_0_61_128 ();
 sg13g2_fill_8 FILLER_0_61_136 ();
 sg13g2_fill_8 FILLER_0_61_144 ();
 sg13g2_fill_8 FILLER_0_61_152 ();
 sg13g2_fill_8 FILLER_0_61_160 ();
 sg13g2_fill_8 FILLER_0_61_168 ();
 sg13g2_fill_8 FILLER_0_61_176 ();
 sg13g2_fill_8 FILLER_0_61_184 ();
 sg13g2_fill_8 FILLER_0_61_192 ();
 sg13g2_fill_8 FILLER_0_61_200 ();
 sg13g2_fill_8 FILLER_0_61_208 ();
 sg13g2_fill_8 FILLER_0_61_216 ();
 sg13g2_fill_2 FILLER_0_61_224 ();
 sg13g2_fill_8 FILLER_0_61_231 ();
 sg13g2_fill_8 FILLER_0_61_239 ();
 sg13g2_fill_4 FILLER_0_61_247 ();
 sg13g2_fill_2 FILLER_0_61_251 ();
 sg13g2_fill_1 FILLER_0_61_253 ();
 sg13g2_fill_2 FILLER_0_61_280 ();
 sg13g2_fill_2 FILLER_0_61_287 ();
 sg13g2_fill_1 FILLER_0_61_289 ();
 sg13g2_fill_2 FILLER_0_61_294 ();
 sg13g2_fill_2 FILLER_0_61_322 ();
 sg13g2_fill_8 FILLER_0_61_350 ();
 sg13g2_fill_4 FILLER_0_61_358 ();
 sg13g2_fill_2 FILLER_0_61_362 ();
 sg13g2_fill_8 FILLER_0_61_369 ();
 sg13g2_fill_8 FILLER_0_61_382 ();
 sg13g2_fill_4 FILLER_0_61_390 ();
 sg13g2_fill_1 FILLER_0_61_394 ();
 sg13g2_fill_2 FILLER_0_61_400 ();
 sg13g2_fill_2 FILLER_0_61_407 ();
 sg13g2_fill_2 FILLER_0_61_415 ();
 sg13g2_fill_4 FILLER_0_61_421 ();
 sg13g2_fill_2 FILLER_0_61_425 ();
 sg13g2_fill_2 FILLER_0_61_432 ();
 sg13g2_fill_4 FILLER_0_61_439 ();
 sg13g2_fill_2 FILLER_0_61_447 ();
 sg13g2_fill_2 FILLER_0_61_455 ();
 sg13g2_fill_1 FILLER_0_61_457 ();
 sg13g2_fill_8 FILLER_0_61_463 ();
 sg13g2_fill_4 FILLER_0_61_471 ();
 sg13g2_fill_1 FILLER_0_61_475 ();
 sg13g2_fill_2 FILLER_0_61_502 ();
 sg13g2_fill_2 FILLER_0_61_509 ();
 sg13g2_fill_2 FILLER_0_61_516 ();
 sg13g2_fill_4 FILLER_0_61_523 ();
 sg13g2_fill_2 FILLER_0_61_533 ();
 sg13g2_fill_2 FILLER_0_61_540 ();
 sg13g2_fill_8 FILLER_0_61_546 ();
 sg13g2_fill_8 FILLER_0_61_554 ();
 sg13g2_fill_8 FILLER_0_61_562 ();
 sg13g2_fill_8 FILLER_0_61_570 ();
 sg13g2_fill_8 FILLER_0_61_578 ();
 sg13g2_fill_8 FILLER_0_61_586 ();
 sg13g2_fill_8 FILLER_0_61_594 ();
 sg13g2_fill_8 FILLER_0_61_602 ();
 sg13g2_fill_8 FILLER_0_61_615 ();
 sg13g2_fill_8 FILLER_0_61_623 ();
 sg13g2_fill_4 FILLER_0_61_657 ();
 sg13g2_fill_1 FILLER_0_61_661 ();
 sg13g2_fill_8 FILLER_0_61_667 ();
 sg13g2_fill_8 FILLER_0_61_680 ();
 sg13g2_fill_8 FILLER_0_61_688 ();
 sg13g2_fill_8 FILLER_0_61_696 ();
 sg13g2_fill_8 FILLER_0_61_704 ();
 sg13g2_fill_8 FILLER_0_61_712 ();
 sg13g2_fill_8 FILLER_0_61_720 ();
 sg13g2_fill_8 FILLER_0_61_728 ();
 sg13g2_fill_4 FILLER_0_61_736 ();
 sg13g2_fill_2 FILLER_0_61_740 ();
 sg13g2_fill_1 FILLER_0_61_742 ();
 sg13g2_fill_8 FILLER_0_61_764 ();
 sg13g2_fill_4 FILLER_0_61_772 ();
 sg13g2_fill_2 FILLER_0_61_780 ();
 sg13g2_fill_8 FILLER_0_61_787 ();
 sg13g2_fill_4 FILLER_0_61_795 ();
 sg13g2_fill_4 FILLER_0_61_804 ();
 sg13g2_fill_8 FILLER_0_61_834 ();
 sg13g2_fill_8 FILLER_0_61_842 ();
 sg13g2_fill_8 FILLER_0_61_850 ();
 sg13g2_fill_4 FILLER_0_61_858 ();
 sg13g2_fill_1 FILLER_0_61_862 ();
 sg13g2_fill_2 FILLER_0_61_868 ();
 sg13g2_fill_1 FILLER_0_61_870 ();
 sg13g2_fill_2 FILLER_0_61_875 ();
 sg13g2_fill_8 FILLER_0_61_882 ();
 sg13g2_fill_8 FILLER_0_61_890 ();
 sg13g2_fill_8 FILLER_0_61_898 ();
 sg13g2_fill_8 FILLER_0_61_906 ();
 sg13g2_fill_8 FILLER_0_61_918 ();
 sg13g2_fill_4 FILLER_0_61_926 ();
 sg13g2_fill_2 FILLER_0_61_930 ();
 sg13g2_fill_4 FILLER_0_61_936 ();
 sg13g2_fill_1 FILLER_0_61_940 ();
 sg13g2_fill_2 FILLER_0_61_945 ();
 sg13g2_fill_2 FILLER_0_61_951 ();
 sg13g2_fill_2 FILLER_0_61_959 ();
 sg13g2_fill_8 FILLER_0_61_964 ();
 sg13g2_fill_4 FILLER_0_61_972 ();
 sg13g2_fill_2 FILLER_0_61_976 ();
 sg13g2_fill_1 FILLER_0_61_978 ();
 sg13g2_fill_8 FILLER_0_61_985 ();
 sg13g2_fill_4 FILLER_0_61_993 ();
 sg13g2_fill_2 FILLER_0_61_997 ();
 sg13g2_fill_4 FILLER_0_61_1005 ();
 sg13g2_fill_8 FILLER_0_61_1017 ();
 sg13g2_fill_1 FILLER_0_61_1025 ();
 sg13g2_fill_4 FILLER_0_61_1031 ();
 sg13g2_fill_1 FILLER_0_61_1035 ();
 sg13g2_fill_2 FILLER_0_61_1041 ();
 sg13g2_fill_8 FILLER_0_61_1050 ();
 sg13g2_fill_8 FILLER_0_61_1058 ();
 sg13g2_fill_4 FILLER_0_61_1066 ();
 sg13g2_fill_1 FILLER_0_61_1070 ();
 sg13g2_fill_2 FILLER_0_61_1076 ();
 sg13g2_fill_2 FILLER_0_61_1082 ();
 sg13g2_fill_1 FILLER_0_61_1084 ();
 sg13g2_fill_2 FILLER_0_61_1090 ();
 sg13g2_fill_2 FILLER_0_61_1097 ();
 sg13g2_fill_2 FILLER_0_61_1105 ();
 sg13g2_fill_4 FILLER_0_61_1112 ();
 sg13g2_fill_8 FILLER_0_61_1121 ();
 sg13g2_fill_2 FILLER_0_61_1129 ();
 sg13g2_fill_8 FILLER_0_61_1136 ();
 sg13g2_fill_8 FILLER_0_61_1144 ();
 sg13g2_fill_8 FILLER_0_61_1152 ();
 sg13g2_fill_8 FILLER_0_61_1160 ();
 sg13g2_fill_2 FILLER_0_61_1168 ();
 sg13g2_fill_1 FILLER_0_61_1170 ();
 sg13g2_fill_8 FILLER_0_61_1175 ();
 sg13g2_fill_8 FILLER_0_61_1183 ();
 sg13g2_fill_8 FILLER_0_61_1191 ();
 sg13g2_fill_1 FILLER_0_61_1199 ();
 sg13g2_fill_4 FILLER_0_61_1205 ();
 sg13g2_fill_2 FILLER_0_61_1214 ();
 sg13g2_fill_8 FILLER_0_61_1223 ();
 sg13g2_fill_1 FILLER_0_61_1231 ();
 sg13g2_fill_8 FILLER_0_61_1237 ();
 sg13g2_fill_4 FILLER_0_61_1245 ();
 sg13g2_fill_2 FILLER_0_61_1249 ();
 sg13g2_fill_1 FILLER_0_61_1251 ();
 sg13g2_fill_2 FILLER_0_61_1257 ();
 sg13g2_fill_4 FILLER_0_61_1264 ();
 sg13g2_fill_2 FILLER_0_61_1272 ();
 sg13g2_fill_2 FILLER_0_61_1279 ();
 sg13g2_fill_4 FILLER_0_61_1286 ();
 sg13g2_fill_2 FILLER_0_61_1290 ();
 sg13g2_fill_1 FILLER_0_61_1296 ();
 sg13g2_fill_8 FILLER_0_62_0 ();
 sg13g2_fill_8 FILLER_0_62_8 ();
 sg13g2_fill_8 FILLER_0_62_16 ();
 sg13g2_fill_8 FILLER_0_62_24 ();
 sg13g2_fill_8 FILLER_0_62_32 ();
 sg13g2_fill_8 FILLER_0_62_40 ();
 sg13g2_fill_8 FILLER_0_62_48 ();
 sg13g2_fill_8 FILLER_0_62_56 ();
 sg13g2_fill_8 FILLER_0_62_64 ();
 sg13g2_fill_8 FILLER_0_62_72 ();
 sg13g2_fill_8 FILLER_0_62_80 ();
 sg13g2_fill_8 FILLER_0_62_88 ();
 sg13g2_fill_8 FILLER_0_62_96 ();
 sg13g2_fill_8 FILLER_0_62_104 ();
 sg13g2_fill_8 FILLER_0_62_112 ();
 sg13g2_fill_8 FILLER_0_62_120 ();
 sg13g2_fill_8 FILLER_0_62_128 ();
 sg13g2_fill_8 FILLER_0_62_136 ();
 sg13g2_fill_8 FILLER_0_62_144 ();
 sg13g2_fill_8 FILLER_0_62_152 ();
 sg13g2_fill_8 FILLER_0_62_160 ();
 sg13g2_fill_8 FILLER_0_62_168 ();
 sg13g2_fill_8 FILLER_0_62_176 ();
 sg13g2_fill_8 FILLER_0_62_184 ();
 sg13g2_fill_8 FILLER_0_62_192 ();
 sg13g2_fill_8 FILLER_0_62_200 ();
 sg13g2_fill_8 FILLER_0_62_208 ();
 sg13g2_fill_8 FILLER_0_62_216 ();
 sg13g2_fill_8 FILLER_0_62_224 ();
 sg13g2_fill_8 FILLER_0_62_232 ();
 sg13g2_fill_8 FILLER_0_62_240 ();
 sg13g2_fill_4 FILLER_0_62_248 ();
 sg13g2_fill_1 FILLER_0_62_252 ();
 sg13g2_fill_8 FILLER_0_62_258 ();
 sg13g2_fill_4 FILLER_0_62_266 ();
 sg13g2_fill_2 FILLER_0_62_270 ();
 sg13g2_fill_8 FILLER_0_62_277 ();
 sg13g2_fill_8 FILLER_0_62_285 ();
 sg13g2_fill_2 FILLER_0_62_293 ();
 sg13g2_fill_1 FILLER_0_62_295 ();
 sg13g2_fill_4 FILLER_0_62_301 ();
 sg13g2_fill_2 FILLER_0_62_305 ();
 sg13g2_fill_4 FILLER_0_62_313 ();
 sg13g2_fill_2 FILLER_0_62_317 ();
 sg13g2_fill_4 FILLER_0_62_331 ();
 sg13g2_fill_2 FILLER_0_62_340 ();
 sg13g2_fill_8 FILLER_0_62_346 ();
 sg13g2_fill_8 FILLER_0_62_380 ();
 sg13g2_fill_4 FILLER_0_62_388 ();
 sg13g2_fill_2 FILLER_0_62_392 ();
 sg13g2_fill_1 FILLER_0_62_394 ();
 sg13g2_fill_2 FILLER_0_62_421 ();
 sg13g2_fill_1 FILLER_0_62_423 ();
 sg13g2_fill_2 FILLER_0_62_429 ();
 sg13g2_fill_2 FILLER_0_62_457 ();
 sg13g2_fill_2 FILLER_0_62_465 ();
 sg13g2_fill_4 FILLER_0_62_472 ();
 sg13g2_fill_2 FILLER_0_62_476 ();
 sg13g2_fill_1 FILLER_0_62_478 ();
 sg13g2_fill_2 FILLER_0_62_505 ();
 sg13g2_fill_4 FILLER_0_62_511 ();
 sg13g2_fill_4 FILLER_0_62_519 ();
 sg13g2_fill_8 FILLER_0_62_549 ();
 sg13g2_fill_8 FILLER_0_62_557 ();
 sg13g2_fill_1 FILLER_0_62_565 ();
 sg13g2_fill_2 FILLER_0_62_570 ();
 sg13g2_fill_8 FILLER_0_62_577 ();
 sg13g2_fill_8 FILLER_0_62_585 ();
 sg13g2_fill_8 FILLER_0_62_593 ();
 sg13g2_fill_2 FILLER_0_62_601 ();
 sg13g2_fill_8 FILLER_0_62_608 ();
 sg13g2_fill_8 FILLER_0_62_616 ();
 sg13g2_fill_4 FILLER_0_62_624 ();
 sg13g2_fill_2 FILLER_0_62_633 ();
 sg13g2_fill_8 FILLER_0_62_639 ();
 sg13g2_fill_2 FILLER_0_62_647 ();
 sg13g2_fill_1 FILLER_0_62_649 ();
 sg13g2_fill_8 FILLER_0_62_654 ();
 sg13g2_fill_8 FILLER_0_62_662 ();
 sg13g2_fill_4 FILLER_0_62_670 ();
 sg13g2_fill_4 FILLER_0_62_683 ();
 sg13g2_fill_2 FILLER_0_62_687 ();
 sg13g2_fill_1 FILLER_0_62_689 ();
 sg13g2_fill_2 FILLER_0_62_695 ();
 sg13g2_fill_2 FILLER_0_62_701 ();
 sg13g2_fill_2 FILLER_0_62_729 ();
 sg13g2_fill_2 FILLER_0_62_736 ();
 sg13g2_fill_8 FILLER_0_62_764 ();
 sg13g2_fill_8 FILLER_0_62_772 ();
 sg13g2_fill_4 FILLER_0_62_780 ();
 sg13g2_fill_2 FILLER_0_62_784 ();
 sg13g2_fill_1 FILLER_0_62_786 ();
 sg13g2_fill_8 FILLER_0_62_792 ();
 sg13g2_fill_8 FILLER_0_62_800 ();
 sg13g2_fill_4 FILLER_0_62_808 ();
 sg13g2_fill_2 FILLER_0_62_817 ();
 sg13g2_fill_8 FILLER_0_62_823 ();
 sg13g2_fill_8 FILLER_0_62_831 ();
 sg13g2_fill_8 FILLER_0_62_839 ();
 sg13g2_fill_8 FILLER_0_62_847 ();
 sg13g2_fill_8 FILLER_0_62_855 ();
 sg13g2_fill_2 FILLER_0_62_868 ();
 sg13g2_fill_2 FILLER_0_62_878 ();
 sg13g2_fill_8 FILLER_0_62_885 ();
 sg13g2_fill_8 FILLER_0_62_893 ();
 sg13g2_fill_8 FILLER_0_62_901 ();
 sg13g2_fill_2 FILLER_0_62_909 ();
 sg13g2_fill_1 FILLER_0_62_911 ();
 sg13g2_fill_4 FILLER_0_62_918 ();
 sg13g2_fill_2 FILLER_0_62_922 ();
 sg13g2_fill_1 FILLER_0_62_924 ();
 sg13g2_fill_4 FILLER_0_62_930 ();
 sg13g2_fill_1 FILLER_0_62_934 ();
 sg13g2_fill_2 FILLER_0_62_945 ();
 sg13g2_fill_8 FILLER_0_62_952 ();
 sg13g2_fill_8 FILLER_0_62_960 ();
 sg13g2_fill_8 FILLER_0_62_968 ();
 sg13g2_fill_4 FILLER_0_62_976 ();
 sg13g2_fill_1 FILLER_0_62_980 ();
 sg13g2_fill_8 FILLER_0_62_986 ();
 sg13g2_fill_4 FILLER_0_62_994 ();
 sg13g2_fill_8 FILLER_0_62_1003 ();
 sg13g2_fill_4 FILLER_0_62_1011 ();
 sg13g2_fill_2 FILLER_0_62_1020 ();
 sg13g2_fill_2 FILLER_0_62_1027 ();
 sg13g2_fill_4 FILLER_0_62_1033 ();
 sg13g2_fill_2 FILLER_0_62_1037 ();
 sg13g2_fill_2 FILLER_0_62_1044 ();
 sg13g2_fill_8 FILLER_0_62_1050 ();
 sg13g2_fill_8 FILLER_0_62_1058 ();
 sg13g2_fill_8 FILLER_0_62_1066 ();
 sg13g2_fill_8 FILLER_0_62_1074 ();
 sg13g2_fill_8 FILLER_0_62_1082 ();
 sg13g2_fill_8 FILLER_0_62_1090 ();
 sg13g2_fill_4 FILLER_0_62_1098 ();
 sg13g2_fill_2 FILLER_0_62_1102 ();
 sg13g2_fill_1 FILLER_0_62_1104 ();
 sg13g2_fill_2 FILLER_0_62_1108 ();
 sg13g2_fill_2 FILLER_0_62_1116 ();
 sg13g2_fill_4 FILLER_0_62_1126 ();
 sg13g2_fill_8 FILLER_0_62_1134 ();
 sg13g2_fill_8 FILLER_0_62_1142 ();
 sg13g2_fill_4 FILLER_0_62_1150 ();
 sg13g2_fill_2 FILLER_0_62_1154 ();
 sg13g2_fill_1 FILLER_0_62_1156 ();
 sg13g2_fill_2 FILLER_0_62_1162 ();
 sg13g2_fill_2 FILLER_0_62_1172 ();
 sg13g2_fill_1 FILLER_0_62_1174 ();
 sg13g2_fill_4 FILLER_0_62_1179 ();
 sg13g2_fill_2 FILLER_0_62_1183 ();
 sg13g2_fill_2 FILLER_0_62_1189 ();
 sg13g2_fill_1 FILLER_0_62_1191 ();
 sg13g2_fill_2 FILLER_0_62_1199 ();
 sg13g2_fill_1 FILLER_0_62_1201 ();
 sg13g2_fill_2 FILLER_0_62_1207 ();
 sg13g2_fill_1 FILLER_0_62_1209 ();
 sg13g2_fill_2 FILLER_0_62_1215 ();
 sg13g2_fill_4 FILLER_0_62_1221 ();
 sg13g2_fill_4 FILLER_0_62_1233 ();
 sg13g2_fill_1 FILLER_0_62_1237 ();
 sg13g2_fill_2 FILLER_0_62_1250 ();
 sg13g2_fill_1 FILLER_0_62_1252 ();
 sg13g2_fill_2 FILLER_0_62_1258 ();
 sg13g2_fill_1 FILLER_0_62_1260 ();
 sg13g2_fill_2 FILLER_0_62_1266 ();
 sg13g2_fill_2 FILLER_0_62_1273 ();
 sg13g2_fill_2 FILLER_0_62_1280 ();
 sg13g2_fill_4 FILLER_0_62_1286 ();
 sg13g2_fill_2 FILLER_0_62_1294 ();
 sg13g2_fill_1 FILLER_0_62_1296 ();
 sg13g2_fill_8 FILLER_0_63_0 ();
 sg13g2_fill_8 FILLER_0_63_8 ();
 sg13g2_fill_8 FILLER_0_63_16 ();
 sg13g2_fill_8 FILLER_0_63_24 ();
 sg13g2_fill_8 FILLER_0_63_32 ();
 sg13g2_fill_8 FILLER_0_63_40 ();
 sg13g2_fill_8 FILLER_0_63_48 ();
 sg13g2_fill_8 FILLER_0_63_56 ();
 sg13g2_fill_8 FILLER_0_63_64 ();
 sg13g2_fill_8 FILLER_0_63_72 ();
 sg13g2_fill_8 FILLER_0_63_80 ();
 sg13g2_fill_8 FILLER_0_63_88 ();
 sg13g2_fill_8 FILLER_0_63_96 ();
 sg13g2_fill_8 FILLER_0_63_104 ();
 sg13g2_fill_8 FILLER_0_63_112 ();
 sg13g2_fill_8 FILLER_0_63_120 ();
 sg13g2_fill_8 FILLER_0_63_128 ();
 sg13g2_fill_8 FILLER_0_63_136 ();
 sg13g2_fill_8 FILLER_0_63_144 ();
 sg13g2_fill_8 FILLER_0_63_152 ();
 sg13g2_fill_8 FILLER_0_63_160 ();
 sg13g2_fill_8 FILLER_0_63_168 ();
 sg13g2_fill_8 FILLER_0_63_176 ();
 sg13g2_fill_8 FILLER_0_63_184 ();
 sg13g2_fill_8 FILLER_0_63_192 ();
 sg13g2_fill_8 FILLER_0_63_200 ();
 sg13g2_fill_8 FILLER_0_63_208 ();
 sg13g2_fill_2 FILLER_0_63_216 ();
 sg13g2_fill_1 FILLER_0_63_218 ();
 sg13g2_fill_2 FILLER_0_63_224 ();
 sg13g2_fill_8 FILLER_0_63_230 ();
 sg13g2_fill_8 FILLER_0_63_238 ();
 sg13g2_fill_8 FILLER_0_63_246 ();
 sg13g2_fill_8 FILLER_0_63_254 ();
 sg13g2_fill_8 FILLER_0_63_262 ();
 sg13g2_fill_8 FILLER_0_63_270 ();
 sg13g2_fill_8 FILLER_0_63_278 ();
 sg13g2_fill_8 FILLER_0_63_286 ();
 sg13g2_fill_8 FILLER_0_63_299 ();
 sg13g2_fill_1 FILLER_0_63_307 ();
 sg13g2_fill_8 FILLER_0_63_313 ();
 sg13g2_fill_8 FILLER_0_63_321 ();
 sg13g2_fill_8 FILLER_0_63_329 ();
 sg13g2_fill_4 FILLER_0_63_337 ();
 sg13g2_fill_8 FILLER_0_63_346 ();
 sg13g2_fill_8 FILLER_0_63_354 ();
 sg13g2_fill_8 FILLER_0_63_362 ();
 sg13g2_fill_8 FILLER_0_63_375 ();
 sg13g2_fill_8 FILLER_0_63_383 ();
 sg13g2_fill_8 FILLER_0_63_391 ();
 sg13g2_fill_8 FILLER_0_63_399 ();
 sg13g2_fill_4 FILLER_0_63_407 ();
 sg13g2_fill_8 FILLER_0_63_416 ();
 sg13g2_fill_8 FILLER_0_63_424 ();
 sg13g2_fill_8 FILLER_0_63_432 ();
 sg13g2_fill_8 FILLER_0_63_440 ();
 sg13g2_fill_4 FILLER_0_63_448 ();
 sg13g2_fill_1 FILLER_0_63_452 ();
 sg13g2_fill_8 FILLER_0_63_458 ();
 sg13g2_fill_8 FILLER_0_63_466 ();
 sg13g2_fill_4 FILLER_0_63_474 ();
 sg13g2_fill_2 FILLER_0_63_478 ();
 sg13g2_fill_1 FILLER_0_63_480 ();
 sg13g2_fill_2 FILLER_0_63_486 ();
 sg13g2_fill_8 FILLER_0_63_492 ();
 sg13g2_fill_8 FILLER_0_63_500 ();
 sg13g2_fill_8 FILLER_0_63_513 ();
 sg13g2_fill_8 FILLER_0_63_521 ();
 sg13g2_fill_8 FILLER_0_63_529 ();
 sg13g2_fill_4 FILLER_0_63_537 ();
 sg13g2_fill_1 FILLER_0_63_541 ();
 sg13g2_fill_2 FILLER_0_63_546 ();
 sg13g2_fill_1 FILLER_0_63_548 ();
 sg13g2_fill_8 FILLER_0_63_554 ();
 sg13g2_fill_1 FILLER_0_63_562 ();
 sg13g2_fill_4 FILLER_0_63_568 ();
 sg13g2_fill_4 FILLER_0_63_577 ();
 sg13g2_fill_1 FILLER_0_63_581 ();
 sg13g2_fill_8 FILLER_0_63_608 ();
 sg13g2_fill_8 FILLER_0_63_616 ();
 sg13g2_fill_4 FILLER_0_63_624 ();
 sg13g2_fill_4 FILLER_0_63_633 ();
 sg13g2_fill_2 FILLER_0_63_637 ();
 sg13g2_fill_1 FILLER_0_63_639 ();
 sg13g2_fill_8 FILLER_0_63_644 ();
 sg13g2_fill_8 FILLER_0_63_652 ();
 sg13g2_fill_8 FILLER_0_63_660 ();
 sg13g2_fill_4 FILLER_0_63_673 ();
 sg13g2_fill_2 FILLER_0_63_677 ();
 sg13g2_fill_1 FILLER_0_63_679 ();
 sg13g2_fill_8 FILLER_0_63_685 ();
 sg13g2_fill_1 FILLER_0_63_693 ();
 sg13g2_fill_2 FILLER_0_63_699 ();
 sg13g2_fill_8 FILLER_0_63_727 ();
 sg13g2_fill_1 FILLER_0_63_735 ();
 sg13g2_fill_4 FILLER_0_63_741 ();
 sg13g2_fill_1 FILLER_0_63_745 ();
 sg13g2_fill_4 FILLER_0_63_750 ();
 sg13g2_fill_1 FILLER_0_63_754 ();
 sg13g2_fill_8 FILLER_0_63_760 ();
 sg13g2_fill_1 FILLER_0_63_768 ();
 sg13g2_fill_2 FILLER_0_63_774 ();
 sg13g2_fill_4 FILLER_0_63_781 ();
 sg13g2_fill_1 FILLER_0_63_785 ();
 sg13g2_fill_4 FILLER_0_63_812 ();
 sg13g2_fill_1 FILLER_0_63_816 ();
 sg13g2_fill_4 FILLER_0_63_838 ();
 sg13g2_fill_2 FILLER_0_63_842 ();
 sg13g2_fill_1 FILLER_0_63_844 ();
 sg13g2_fill_8 FILLER_0_63_850 ();
 sg13g2_fill_8 FILLER_0_63_884 ();
 sg13g2_fill_4 FILLER_0_63_892 ();
 sg13g2_fill_2 FILLER_0_63_896 ();
 sg13g2_fill_8 FILLER_0_63_903 ();
 sg13g2_fill_4 FILLER_0_63_911 ();
 sg13g2_fill_1 FILLER_0_63_915 ();
 sg13g2_fill_2 FILLER_0_63_920 ();
 sg13g2_fill_1 FILLER_0_63_922 ();
 sg13g2_fill_8 FILLER_0_63_927 ();
 sg13g2_fill_2 FILLER_0_63_940 ();
 sg13g2_fill_8 FILLER_0_63_946 ();
 sg13g2_fill_2 FILLER_0_63_959 ();
 sg13g2_fill_8 FILLER_0_63_967 ();
 sg13g2_fill_2 FILLER_0_63_979 ();
 sg13g2_fill_2 FILLER_0_63_993 ();
 sg13g2_fill_2 FILLER_0_63_1001 ();
 sg13g2_fill_2 FILLER_0_63_1008 ();
 sg13g2_fill_2 FILLER_0_63_1015 ();
 sg13g2_fill_4 FILLER_0_63_1022 ();
 sg13g2_fill_2 FILLER_0_63_1026 ();
 sg13g2_fill_1 FILLER_0_63_1028 ();
 sg13g2_fill_4 FILLER_0_63_1034 ();
 sg13g2_fill_1 FILLER_0_63_1038 ();
 sg13g2_fill_2 FILLER_0_63_1043 ();
 sg13g2_fill_2 FILLER_0_63_1050 ();
 sg13g2_fill_8 FILLER_0_63_1057 ();
 sg13g2_fill_8 FILLER_0_63_1065 ();
 sg13g2_fill_8 FILLER_0_63_1073 ();
 sg13g2_fill_2 FILLER_0_63_1086 ();
 sg13g2_fill_8 FILLER_0_63_1092 ();
 sg13g2_fill_4 FILLER_0_63_1100 ();
 sg13g2_fill_2 FILLER_0_63_1104 ();
 sg13g2_fill_2 FILLER_0_63_1111 ();
 sg13g2_fill_8 FILLER_0_63_1118 ();
 sg13g2_fill_4 FILLER_0_63_1126 ();
 sg13g2_fill_2 FILLER_0_63_1130 ();
 sg13g2_fill_4 FILLER_0_63_1138 ();
 sg13g2_fill_2 FILLER_0_63_1146 ();
 sg13g2_fill_2 FILLER_0_63_1152 ();
 sg13g2_fill_1 FILLER_0_63_1154 ();
 sg13g2_fill_2 FILLER_0_63_1160 ();
 sg13g2_fill_2 FILLER_0_63_1170 ();
 sg13g2_fill_1 FILLER_0_63_1172 ();
 sg13g2_fill_2 FILLER_0_63_1177 ();
 sg13g2_fill_2 FILLER_0_63_1185 ();
 sg13g2_fill_4 FILLER_0_63_1192 ();
 sg13g2_fill_1 FILLER_0_63_1196 ();
 sg13g2_fill_8 FILLER_0_63_1203 ();
 sg13g2_fill_8 FILLER_0_63_1214 ();
 sg13g2_fill_8 FILLER_0_63_1222 ();
 sg13g2_fill_4 FILLER_0_63_1230 ();
 sg13g2_fill_2 FILLER_0_63_1234 ();
 sg13g2_fill_2 FILLER_0_63_1241 ();
 sg13g2_fill_2 FILLER_0_63_1249 ();
 sg13g2_fill_2 FILLER_0_63_1256 ();
 sg13g2_fill_2 FILLER_0_63_1262 ();
 sg13g2_fill_1 FILLER_0_63_1264 ();
 sg13g2_fill_2 FILLER_0_63_1270 ();
 sg13g2_fill_4 FILLER_0_63_1277 ();
 sg13g2_fill_2 FILLER_0_63_1286 ();
 sg13g2_fill_4 FILLER_0_63_1293 ();
 sg13g2_fill_8 FILLER_0_64_0 ();
 sg13g2_fill_8 FILLER_0_64_8 ();
 sg13g2_fill_8 FILLER_0_64_16 ();
 sg13g2_fill_8 FILLER_0_64_24 ();
 sg13g2_fill_8 FILLER_0_64_32 ();
 sg13g2_fill_8 FILLER_0_64_40 ();
 sg13g2_fill_8 FILLER_0_64_48 ();
 sg13g2_fill_8 FILLER_0_64_56 ();
 sg13g2_fill_8 FILLER_0_64_64 ();
 sg13g2_fill_8 FILLER_0_64_72 ();
 sg13g2_fill_8 FILLER_0_64_80 ();
 sg13g2_fill_8 FILLER_0_64_88 ();
 sg13g2_fill_8 FILLER_0_64_96 ();
 sg13g2_fill_8 FILLER_0_64_104 ();
 sg13g2_fill_8 FILLER_0_64_112 ();
 sg13g2_fill_8 FILLER_0_64_120 ();
 sg13g2_fill_8 FILLER_0_64_128 ();
 sg13g2_fill_8 FILLER_0_64_136 ();
 sg13g2_fill_8 FILLER_0_64_144 ();
 sg13g2_fill_8 FILLER_0_64_152 ();
 sg13g2_fill_8 FILLER_0_64_160 ();
 sg13g2_fill_8 FILLER_0_64_168 ();
 sg13g2_fill_8 FILLER_0_64_176 ();
 sg13g2_fill_8 FILLER_0_64_184 ();
 sg13g2_fill_8 FILLER_0_64_192 ();
 sg13g2_fill_8 FILLER_0_64_200 ();
 sg13g2_fill_4 FILLER_0_64_208 ();
 sg13g2_fill_2 FILLER_0_64_212 ();
 sg13g2_fill_2 FILLER_0_64_240 ();
 sg13g2_fill_1 FILLER_0_64_242 ();
 sg13g2_fill_4 FILLER_0_64_247 ();
 sg13g2_fill_4 FILLER_0_64_257 ();
 sg13g2_fill_2 FILLER_0_64_261 ();
 sg13g2_fill_1 FILLER_0_64_263 ();
 sg13g2_fill_2 FILLER_0_64_269 ();
 sg13g2_fill_2 FILLER_0_64_277 ();
 sg13g2_fill_8 FILLER_0_64_285 ();
 sg13g2_fill_8 FILLER_0_64_293 ();
 sg13g2_fill_4 FILLER_0_64_301 ();
 sg13g2_fill_2 FILLER_0_64_305 ();
 sg13g2_fill_1 FILLER_0_64_307 ();
 sg13g2_fill_8 FILLER_0_64_314 ();
 sg13g2_fill_2 FILLER_0_64_322 ();
 sg13g2_fill_2 FILLER_0_64_332 ();
 sg13g2_fill_2 FILLER_0_64_344 ();
 sg13g2_fill_8 FILLER_0_64_351 ();
 sg13g2_fill_2 FILLER_0_64_359 ();
 sg13g2_fill_4 FILLER_0_64_368 ();
 sg13g2_fill_1 FILLER_0_64_372 ();
 sg13g2_fill_8 FILLER_0_64_378 ();
 sg13g2_fill_8 FILLER_0_64_386 ();
 sg13g2_fill_8 FILLER_0_64_394 ();
 sg13g2_fill_8 FILLER_0_64_402 ();
 sg13g2_fill_8 FILLER_0_64_410 ();
 sg13g2_fill_4 FILLER_0_64_418 ();
 sg13g2_fill_1 FILLER_0_64_422 ();
 sg13g2_fill_8 FILLER_0_64_428 ();
 sg13g2_fill_1 FILLER_0_64_436 ();
 sg13g2_fill_8 FILLER_0_64_443 ();
 sg13g2_fill_8 FILLER_0_64_451 ();
 sg13g2_fill_8 FILLER_0_64_459 ();
 sg13g2_fill_8 FILLER_0_64_467 ();
 sg13g2_fill_8 FILLER_0_64_475 ();
 sg13g2_fill_8 FILLER_0_64_483 ();
 sg13g2_fill_8 FILLER_0_64_491 ();
 sg13g2_fill_8 FILLER_0_64_499 ();
 sg13g2_fill_8 FILLER_0_64_507 ();
 sg13g2_fill_8 FILLER_0_64_515 ();
 sg13g2_fill_8 FILLER_0_64_523 ();
 sg13g2_fill_8 FILLER_0_64_531 ();
 sg13g2_fill_2 FILLER_0_64_546 ();
 sg13g2_fill_2 FILLER_0_64_574 ();
 sg13g2_fill_4 FILLER_0_64_580 ();
 sg13g2_fill_8 FILLER_0_64_605 ();
 sg13g2_fill_8 FILLER_0_64_613 ();
 sg13g2_fill_2 FILLER_0_64_621 ();
 sg13g2_fill_8 FILLER_0_64_649 ();
 sg13g2_fill_2 FILLER_0_64_657 ();
 sg13g2_fill_8 FILLER_0_64_685 ();
 sg13g2_fill_8 FILLER_0_64_693 ();
 sg13g2_fill_8 FILLER_0_64_701 ();
 sg13g2_fill_2 FILLER_0_64_709 ();
 sg13g2_fill_4 FILLER_0_64_716 ();
 sg13g2_fill_2 FILLER_0_64_720 ();
 sg13g2_fill_1 FILLER_0_64_722 ();
 sg13g2_fill_8 FILLER_0_64_733 ();
 sg13g2_fill_4 FILLER_0_64_741 ();
 sg13g2_fill_1 FILLER_0_64_745 ();
 sg13g2_fill_8 FILLER_0_64_751 ();
 sg13g2_fill_1 FILLER_0_64_759 ();
 sg13g2_fill_2 FILLER_0_64_765 ();
 sg13g2_fill_2 FILLER_0_64_793 ();
 sg13g2_fill_2 FILLER_0_64_799 ();
 sg13g2_fill_4 FILLER_0_64_806 ();
 sg13g2_fill_2 FILLER_0_64_836 ();
 sg13g2_fill_8 FILLER_0_64_843 ();
 sg13g2_fill_8 FILLER_0_64_851 ();
 sg13g2_fill_4 FILLER_0_64_859 ();
 sg13g2_fill_2 FILLER_0_64_863 ();
 sg13g2_fill_1 FILLER_0_64_865 ();
 sg13g2_fill_8 FILLER_0_64_871 ();
 sg13g2_fill_8 FILLER_0_64_879 ();
 sg13g2_fill_8 FILLER_0_64_887 ();
 sg13g2_fill_2 FILLER_0_64_895 ();
 sg13g2_fill_2 FILLER_0_64_901 ();
 sg13g2_fill_4 FILLER_0_64_907 ();
 sg13g2_fill_1 FILLER_0_64_911 ();
 sg13g2_fill_8 FILLER_0_64_917 ();
 sg13g2_fill_8 FILLER_0_64_925 ();
 sg13g2_fill_8 FILLER_0_64_933 ();
 sg13g2_fill_4 FILLER_0_64_941 ();
 sg13g2_fill_8 FILLER_0_64_951 ();
 sg13g2_fill_1 FILLER_0_64_959 ();
 sg13g2_fill_2 FILLER_0_64_964 ();
 sg13g2_fill_4 FILLER_0_64_971 ();
 sg13g2_fill_8 FILLER_0_64_980 ();
 sg13g2_fill_8 FILLER_0_64_988 ();
 sg13g2_fill_1 FILLER_0_64_996 ();
 sg13g2_fill_2 FILLER_0_64_1002 ();
 sg13g2_fill_4 FILLER_0_64_1008 ();
 sg13g2_fill_2 FILLER_0_64_1017 ();
 sg13g2_fill_1 FILLER_0_64_1019 ();
 sg13g2_fill_2 FILLER_0_64_1024 ();
 sg13g2_fill_2 FILLER_0_64_1033 ();
 sg13g2_fill_2 FILLER_0_64_1041 ();
 sg13g2_fill_2 FILLER_0_64_1048 ();
 sg13g2_fill_8 FILLER_0_64_1056 ();
 sg13g2_fill_2 FILLER_0_64_1064 ();
 sg13g2_fill_1 FILLER_0_64_1066 ();
 sg13g2_fill_8 FILLER_0_64_1072 ();
 sg13g2_fill_4 FILLER_0_64_1080 ();
 sg13g2_fill_1 FILLER_0_64_1084 ();
 sg13g2_fill_8 FILLER_0_64_1089 ();
 sg13g2_fill_8 FILLER_0_64_1097 ();
 sg13g2_fill_4 FILLER_0_64_1105 ();
 sg13g2_fill_2 FILLER_0_64_1113 ();
 sg13g2_fill_1 FILLER_0_64_1115 ();
 sg13g2_fill_8 FILLER_0_64_1120 ();
 sg13g2_fill_1 FILLER_0_64_1128 ();
 sg13g2_fill_2 FILLER_0_64_1137 ();
 sg13g2_fill_8 FILLER_0_64_1144 ();
 sg13g2_fill_8 FILLER_0_64_1152 ();
 sg13g2_fill_8 FILLER_0_64_1160 ();
 sg13g2_fill_8 FILLER_0_64_1168 ();
 sg13g2_fill_4 FILLER_0_64_1176 ();
 sg13g2_fill_2 FILLER_0_64_1180 ();
 sg13g2_fill_2 FILLER_0_64_1189 ();
 sg13g2_fill_2 FILLER_0_64_1197 ();
 sg13g2_fill_1 FILLER_0_64_1199 ();
 sg13g2_fill_2 FILLER_0_64_1204 ();
 sg13g2_fill_8 FILLER_0_64_1211 ();
 sg13g2_fill_8 FILLER_0_64_1219 ();
 sg13g2_fill_8 FILLER_0_64_1227 ();
 sg13g2_fill_1 FILLER_0_64_1235 ();
 sg13g2_fill_8 FILLER_0_64_1240 ();
 sg13g2_fill_8 FILLER_0_64_1248 ();
 sg13g2_fill_2 FILLER_0_64_1256 ();
 sg13g2_fill_1 FILLER_0_64_1258 ();
 sg13g2_fill_8 FILLER_0_64_1263 ();
 sg13g2_fill_8 FILLER_0_64_1271 ();
 sg13g2_fill_2 FILLER_0_64_1284 ();
 sg13g2_fill_2 FILLER_0_64_1290 ();
 sg13g2_fill_1 FILLER_0_64_1296 ();
 sg13g2_fill_8 FILLER_0_65_0 ();
 sg13g2_fill_8 FILLER_0_65_8 ();
 sg13g2_fill_8 FILLER_0_65_16 ();
 sg13g2_fill_8 FILLER_0_65_24 ();
 sg13g2_fill_8 FILLER_0_65_32 ();
 sg13g2_fill_8 FILLER_0_65_40 ();
 sg13g2_fill_8 FILLER_0_65_48 ();
 sg13g2_fill_8 FILLER_0_65_56 ();
 sg13g2_fill_8 FILLER_0_65_64 ();
 sg13g2_fill_8 FILLER_0_65_72 ();
 sg13g2_fill_8 FILLER_0_65_80 ();
 sg13g2_fill_8 FILLER_0_65_88 ();
 sg13g2_fill_8 FILLER_0_65_96 ();
 sg13g2_fill_8 FILLER_0_65_104 ();
 sg13g2_fill_8 FILLER_0_65_112 ();
 sg13g2_fill_8 FILLER_0_65_120 ();
 sg13g2_fill_8 FILLER_0_65_128 ();
 sg13g2_fill_8 FILLER_0_65_136 ();
 sg13g2_fill_8 FILLER_0_65_144 ();
 sg13g2_fill_8 FILLER_0_65_152 ();
 sg13g2_fill_8 FILLER_0_65_160 ();
 sg13g2_fill_8 FILLER_0_65_168 ();
 sg13g2_fill_8 FILLER_0_65_176 ();
 sg13g2_fill_8 FILLER_0_65_184 ();
 sg13g2_fill_8 FILLER_0_65_192 ();
 sg13g2_fill_8 FILLER_0_65_200 ();
 sg13g2_fill_8 FILLER_0_65_208 ();
 sg13g2_fill_8 FILLER_0_65_216 ();
 sg13g2_fill_4 FILLER_0_65_224 ();
 sg13g2_fill_2 FILLER_0_65_228 ();
 sg13g2_fill_1 FILLER_0_65_230 ();
 sg13g2_fill_2 FILLER_0_65_257 ();
 sg13g2_fill_2 FILLER_0_65_285 ();
 sg13g2_fill_4 FILLER_0_65_291 ();
 sg13g2_fill_2 FILLER_0_65_300 ();
 sg13g2_fill_4 FILLER_0_65_306 ();
 sg13g2_fill_1 FILLER_0_65_310 ();
 sg13g2_fill_2 FILLER_0_65_337 ();
 sg13g2_fill_8 FILLER_0_65_343 ();
 sg13g2_fill_4 FILLER_0_65_351 ();
 sg13g2_fill_2 FILLER_0_65_363 ();
 sg13g2_fill_2 FILLER_0_65_370 ();
 sg13g2_fill_2 FILLER_0_65_376 ();
 sg13g2_fill_8 FILLER_0_65_383 ();
 sg13g2_fill_4 FILLER_0_65_391 ();
 sg13g2_fill_2 FILLER_0_65_395 ();
 sg13g2_fill_1 FILLER_0_65_397 ();
 sg13g2_fill_4 FILLER_0_65_403 ();
 sg13g2_fill_2 FILLER_0_65_412 ();
 sg13g2_fill_8 FILLER_0_65_424 ();
 sg13g2_fill_8 FILLER_0_65_432 ();
 sg13g2_fill_8 FILLER_0_65_440 ();
 sg13g2_fill_4 FILLER_0_65_448 ();
 sg13g2_fill_1 FILLER_0_65_452 ();
 sg13g2_fill_2 FILLER_0_65_458 ();
 sg13g2_fill_1 FILLER_0_65_460 ();
 sg13g2_fill_8 FILLER_0_65_465 ();
 sg13g2_fill_8 FILLER_0_65_473 ();
 sg13g2_fill_2 FILLER_0_65_481 ();
 sg13g2_fill_2 FILLER_0_65_487 ();
 sg13g2_fill_8 FILLER_0_65_515 ();
 sg13g2_fill_1 FILLER_0_65_523 ();
 sg13g2_fill_8 FILLER_0_65_529 ();
 sg13g2_fill_8 FILLER_0_65_537 ();
 sg13g2_fill_1 FILLER_0_65_545 ();
 sg13g2_fill_8 FILLER_0_65_554 ();
 sg13g2_fill_2 FILLER_0_65_562 ();
 sg13g2_fill_8 FILLER_0_65_568 ();
 sg13g2_fill_2 FILLER_0_65_576 ();
 sg13g2_fill_1 FILLER_0_65_578 ();
 sg13g2_fill_4 FILLER_0_65_589 ();
 sg13g2_fill_1 FILLER_0_65_593 ();
 sg13g2_fill_2 FILLER_0_65_599 ();
 sg13g2_fill_8 FILLER_0_65_605 ();
 sg13g2_fill_8 FILLER_0_65_613 ();
 sg13g2_fill_8 FILLER_0_65_621 ();
 sg13g2_fill_8 FILLER_0_65_629 ();
 sg13g2_fill_8 FILLER_0_65_637 ();
 sg13g2_fill_2 FILLER_0_65_666 ();
 sg13g2_fill_2 FILLER_0_65_672 ();
 sg13g2_fill_1 FILLER_0_65_674 ();
 sg13g2_fill_8 FILLER_0_65_679 ();
 sg13g2_fill_8 FILLER_0_65_687 ();
 sg13g2_fill_8 FILLER_0_65_695 ();
 sg13g2_fill_8 FILLER_0_65_703 ();
 sg13g2_fill_8 FILLER_0_65_715 ();
 sg13g2_fill_8 FILLER_0_65_723 ();
 sg13g2_fill_4 FILLER_0_65_731 ();
 sg13g2_fill_2 FILLER_0_65_740 ();
 sg13g2_fill_1 FILLER_0_65_742 ();
 sg13g2_fill_8 FILLER_0_65_748 ();
 sg13g2_fill_8 FILLER_0_65_756 ();
 sg13g2_fill_8 FILLER_0_65_764 ();
 sg13g2_fill_4 FILLER_0_65_772 ();
 sg13g2_fill_2 FILLER_0_65_776 ();
 sg13g2_fill_8 FILLER_0_65_782 ();
 sg13g2_fill_4 FILLER_0_65_790 ();
 sg13g2_fill_2 FILLER_0_65_794 ();
 sg13g2_fill_2 FILLER_0_65_806 ();
 sg13g2_fill_4 FILLER_0_65_812 ();
 sg13g2_fill_2 FILLER_0_65_816 ();
 sg13g2_fill_1 FILLER_0_65_818 ();
 sg13g2_fill_2 FILLER_0_65_824 ();
 sg13g2_fill_2 FILLER_0_65_836 ();
 sg13g2_fill_8 FILLER_0_65_842 ();
 sg13g2_fill_8 FILLER_0_65_850 ();
 sg13g2_fill_4 FILLER_0_65_858 ();
 sg13g2_fill_1 FILLER_0_65_862 ();
 sg13g2_fill_2 FILLER_0_65_871 ();
 sg13g2_fill_1 FILLER_0_65_873 ();
 sg13g2_fill_8 FILLER_0_65_882 ();
 sg13g2_fill_8 FILLER_0_65_890 ();
 sg13g2_fill_4 FILLER_0_65_898 ();
 sg13g2_fill_2 FILLER_0_65_902 ();
 sg13g2_fill_2 FILLER_0_65_909 ();
 sg13g2_fill_4 FILLER_0_65_921 ();
 sg13g2_fill_2 FILLER_0_65_925 ();
 sg13g2_fill_1 FILLER_0_65_927 ();
 sg13g2_fill_2 FILLER_0_65_933 ();
 sg13g2_fill_2 FILLER_0_65_940 ();
 sg13g2_fill_1 FILLER_0_65_942 ();
 sg13g2_fill_2 FILLER_0_65_947 ();
 sg13g2_fill_2 FILLER_0_65_954 ();
 sg13g2_fill_8 FILLER_0_65_963 ();
 sg13g2_fill_8 FILLER_0_65_976 ();
 sg13g2_fill_8 FILLER_0_65_984 ();
 sg13g2_fill_8 FILLER_0_65_992 ();
 sg13g2_fill_1 FILLER_0_65_1000 ();
 sg13g2_fill_4 FILLER_0_65_1008 ();
 sg13g2_fill_1 FILLER_0_65_1012 ();
 sg13g2_fill_2 FILLER_0_65_1018 ();
 sg13g2_fill_4 FILLER_0_65_1025 ();
 sg13g2_fill_1 FILLER_0_65_1029 ();
 sg13g2_fill_2 FILLER_0_65_1034 ();
 sg13g2_fill_4 FILLER_0_65_1041 ();
 sg13g2_fill_2 FILLER_0_65_1045 ();
 sg13g2_fill_2 FILLER_0_65_1054 ();
 sg13g2_fill_2 FILLER_0_65_1060 ();
 sg13g2_fill_8 FILLER_0_65_1068 ();
 sg13g2_fill_8 FILLER_0_65_1076 ();
 sg13g2_fill_2 FILLER_0_65_1084 ();
 sg13g2_fill_8 FILLER_0_65_1091 ();
 sg13g2_fill_8 FILLER_0_65_1099 ();
 sg13g2_fill_4 FILLER_0_65_1107 ();
 sg13g2_fill_2 FILLER_0_65_1118 ();
 sg13g2_fill_8 FILLER_0_65_1124 ();
 sg13g2_fill_8 FILLER_0_65_1132 ();
 sg13g2_fill_8 FILLER_0_65_1140 ();
 sg13g2_fill_8 FILLER_0_65_1148 ();
 sg13g2_fill_8 FILLER_0_65_1156 ();
 sg13g2_fill_4 FILLER_0_65_1164 ();
 sg13g2_fill_2 FILLER_0_65_1168 ();
 sg13g2_fill_4 FILLER_0_65_1178 ();
 sg13g2_fill_2 FILLER_0_65_1182 ();
 sg13g2_fill_1 FILLER_0_65_1184 ();
 sg13g2_fill_2 FILLER_0_65_1189 ();
 sg13g2_fill_8 FILLER_0_65_1195 ();
 sg13g2_fill_1 FILLER_0_65_1203 ();
 sg13g2_fill_2 FILLER_0_65_1209 ();
 sg13g2_fill_8 FILLER_0_65_1214 ();
 sg13g2_fill_2 FILLER_0_65_1222 ();
 sg13g2_fill_1 FILLER_0_65_1224 ();
 sg13g2_fill_8 FILLER_0_65_1230 ();
 sg13g2_fill_8 FILLER_0_65_1238 ();
 sg13g2_fill_8 FILLER_0_65_1246 ();
 sg13g2_fill_4 FILLER_0_65_1260 ();
 sg13g2_fill_2 FILLER_0_65_1268 ();
 sg13g2_fill_8 FILLER_0_65_1277 ();
 sg13g2_fill_2 FILLER_0_65_1289 ();
 sg13g2_fill_2 FILLER_0_65_1295 ();
 sg13g2_fill_8 FILLER_0_66_0 ();
 sg13g2_fill_8 FILLER_0_66_8 ();
 sg13g2_fill_8 FILLER_0_66_16 ();
 sg13g2_fill_8 FILLER_0_66_24 ();
 sg13g2_fill_8 FILLER_0_66_32 ();
 sg13g2_fill_8 FILLER_0_66_40 ();
 sg13g2_fill_8 FILLER_0_66_48 ();
 sg13g2_fill_8 FILLER_0_66_56 ();
 sg13g2_fill_8 FILLER_0_66_64 ();
 sg13g2_fill_8 FILLER_0_66_72 ();
 sg13g2_fill_8 FILLER_0_66_80 ();
 sg13g2_fill_8 FILLER_0_66_88 ();
 sg13g2_fill_8 FILLER_0_66_96 ();
 sg13g2_fill_8 FILLER_0_66_104 ();
 sg13g2_fill_8 FILLER_0_66_112 ();
 sg13g2_fill_8 FILLER_0_66_120 ();
 sg13g2_fill_8 FILLER_0_66_128 ();
 sg13g2_fill_8 FILLER_0_66_136 ();
 sg13g2_fill_4 FILLER_0_66_144 ();
 sg13g2_fill_2 FILLER_0_66_148 ();
 sg13g2_fill_1 FILLER_0_66_150 ();
 sg13g2_fill_8 FILLER_0_66_155 ();
 sg13g2_fill_8 FILLER_0_66_163 ();
 sg13g2_fill_8 FILLER_0_66_171 ();
 sg13g2_fill_8 FILLER_0_66_179 ();
 sg13g2_fill_8 FILLER_0_66_187 ();
 sg13g2_fill_8 FILLER_0_66_195 ();
 sg13g2_fill_8 FILLER_0_66_203 ();
 sg13g2_fill_8 FILLER_0_66_211 ();
 sg13g2_fill_8 FILLER_0_66_219 ();
 sg13g2_fill_4 FILLER_0_66_227 ();
 sg13g2_fill_2 FILLER_0_66_231 ();
 sg13g2_fill_2 FILLER_0_66_238 ();
 sg13g2_fill_4 FILLER_0_66_245 ();
 sg13g2_fill_2 FILLER_0_66_249 ();
 sg13g2_fill_1 FILLER_0_66_251 ();
 sg13g2_fill_2 FILLER_0_66_258 ();
 sg13g2_fill_8 FILLER_0_66_265 ();
 sg13g2_fill_1 FILLER_0_66_273 ();
 sg13g2_fill_8 FILLER_0_66_279 ();
 sg13g2_fill_2 FILLER_0_66_292 ();
 sg13g2_fill_2 FILLER_0_66_299 ();
 sg13g2_fill_8 FILLER_0_66_307 ();
 sg13g2_fill_8 FILLER_0_66_315 ();
 sg13g2_fill_8 FILLER_0_66_323 ();
 sg13g2_fill_1 FILLER_0_66_331 ();
 sg13g2_fill_2 FILLER_0_66_337 ();
 sg13g2_fill_1 FILLER_0_66_339 ();
 sg13g2_fill_2 FILLER_0_66_366 ();
 sg13g2_fill_2 FILLER_0_66_373 ();
 sg13g2_fill_8 FILLER_0_66_380 ();
 sg13g2_fill_8 FILLER_0_66_388 ();
 sg13g2_fill_2 FILLER_0_66_396 ();
 sg13g2_fill_4 FILLER_0_66_402 ();
 sg13g2_fill_2 FILLER_0_66_432 ();
 sg13g2_fill_4 FILLER_0_66_438 ();
 sg13g2_fill_2 FILLER_0_66_447 ();
 sg13g2_fill_2 FILLER_0_66_475 ();
 sg13g2_fill_2 FILLER_0_66_482 ();
 sg13g2_fill_4 FILLER_0_66_489 ();
 sg13g2_fill_2 FILLER_0_66_519 ();
 sg13g2_fill_8 FILLER_0_66_542 ();
 sg13g2_fill_8 FILLER_0_66_550 ();
 sg13g2_fill_8 FILLER_0_66_558 ();
 sg13g2_fill_8 FILLER_0_66_566 ();
 sg13g2_fill_8 FILLER_0_66_574 ();
 sg13g2_fill_4 FILLER_0_66_582 ();
 sg13g2_fill_2 FILLER_0_66_591 ();
 sg13g2_fill_2 FILLER_0_66_598 ();
 sg13g2_fill_8 FILLER_0_66_605 ();
 sg13g2_fill_8 FILLER_0_66_613 ();
 sg13g2_fill_2 FILLER_0_66_621 ();
 sg13g2_fill_2 FILLER_0_66_628 ();
 sg13g2_fill_8 FILLER_0_66_656 ();
 sg13g2_fill_1 FILLER_0_66_664 ();
 sg13g2_fill_8 FILLER_0_66_686 ();
 sg13g2_fill_8 FILLER_0_66_694 ();
 sg13g2_fill_8 FILLER_0_66_702 ();
 sg13g2_fill_8 FILLER_0_66_710 ();
 sg13g2_fill_8 FILLER_0_66_718 ();
 sg13g2_fill_4 FILLER_0_66_726 ();
 sg13g2_fill_2 FILLER_0_66_730 ();
 sg13g2_fill_1 FILLER_0_66_732 ();
 sg13g2_fill_2 FILLER_0_66_759 ();
 sg13g2_fill_8 FILLER_0_66_765 ();
 sg13g2_fill_8 FILLER_0_66_773 ();
 sg13g2_fill_8 FILLER_0_66_781 ();
 sg13g2_fill_8 FILLER_0_66_789 ();
 sg13g2_fill_8 FILLER_0_66_797 ();
 sg13g2_fill_8 FILLER_0_66_810 ();
 sg13g2_fill_8 FILLER_0_66_822 ();
 sg13g2_fill_8 FILLER_0_66_830 ();
 sg13g2_fill_8 FILLER_0_66_838 ();
 sg13g2_fill_8 FILLER_0_66_846 ();
 sg13g2_fill_8 FILLER_0_66_854 ();
 sg13g2_fill_8 FILLER_0_66_862 ();
 sg13g2_fill_8 FILLER_0_66_870 ();
 sg13g2_fill_8 FILLER_0_66_878 ();
 sg13g2_fill_8 FILLER_0_66_886 ();
 sg13g2_fill_4 FILLER_0_66_894 ();
 sg13g2_fill_8 FILLER_0_66_902 ();
 sg13g2_fill_4 FILLER_0_66_910 ();
 sg13g2_fill_1 FILLER_0_66_914 ();
 sg13g2_fill_8 FILLER_0_66_919 ();
 sg13g2_fill_1 FILLER_0_66_927 ();
 sg13g2_fill_2 FILLER_0_66_934 ();
 sg13g2_fill_2 FILLER_0_66_940 ();
 sg13g2_fill_8 FILLER_0_66_947 ();
 sg13g2_fill_8 FILLER_0_66_955 ();
 sg13g2_fill_8 FILLER_0_66_963 ();
 sg13g2_fill_8 FILLER_0_66_971 ();
 sg13g2_fill_4 FILLER_0_66_979 ();
 sg13g2_fill_1 FILLER_0_66_983 ();
 sg13g2_fill_8 FILLER_0_66_989 ();
 sg13g2_fill_8 FILLER_0_66_997 ();
 sg13g2_fill_4 FILLER_0_66_1005 ();
 sg13g2_fill_8 FILLER_0_66_1013 ();
 sg13g2_fill_8 FILLER_0_66_1021 ();
 sg13g2_fill_8 FILLER_0_66_1029 ();
 sg13g2_fill_8 FILLER_0_66_1037 ();
 sg13g2_fill_4 FILLER_0_66_1049 ();
 sg13g2_fill_8 FILLER_0_66_1058 ();
 sg13g2_fill_8 FILLER_0_66_1066 ();
 sg13g2_fill_8 FILLER_0_66_1074 ();
 sg13g2_fill_8 FILLER_0_66_1082 ();
 sg13g2_fill_8 FILLER_0_66_1090 ();
 sg13g2_fill_8 FILLER_0_66_1098 ();
 sg13g2_fill_8 FILLER_0_66_1106 ();
 sg13g2_fill_4 FILLER_0_66_1114 ();
 sg13g2_fill_2 FILLER_0_66_1118 ();
 sg13g2_fill_8 FILLER_0_66_1125 ();
 sg13g2_fill_1 FILLER_0_66_1133 ();
 sg13g2_fill_8 FILLER_0_66_1137 ();
 sg13g2_fill_1 FILLER_0_66_1145 ();
 sg13g2_fill_4 FILLER_0_66_1150 ();
 sg13g2_fill_8 FILLER_0_66_1158 ();
 sg13g2_fill_8 FILLER_0_66_1166 ();
 sg13g2_fill_8 FILLER_0_66_1174 ();
 sg13g2_fill_2 FILLER_0_66_1188 ();
 sg13g2_fill_8 FILLER_0_66_1193 ();
 sg13g2_fill_8 FILLER_0_66_1201 ();
 sg13g2_fill_8 FILLER_0_66_1209 ();
 sg13g2_fill_4 FILLER_0_66_1217 ();
 sg13g2_fill_2 FILLER_0_66_1221 ();
 sg13g2_fill_4 FILLER_0_66_1227 ();
 sg13g2_fill_2 FILLER_0_66_1235 ();
 sg13g2_fill_8 FILLER_0_66_1242 ();
 sg13g2_fill_8 FILLER_0_66_1250 ();
 sg13g2_fill_2 FILLER_0_66_1258 ();
 sg13g2_fill_8 FILLER_0_66_1263 ();
 sg13g2_fill_8 FILLER_0_66_1275 ();
 sg13g2_fill_2 FILLER_0_66_1283 ();
 sg13g2_fill_2 FILLER_0_66_1290 ();
 sg13g2_fill_1 FILLER_0_66_1296 ();
 sg13g2_fill_8 FILLER_0_67_0 ();
 sg13g2_fill_8 FILLER_0_67_8 ();
 sg13g2_fill_8 FILLER_0_67_16 ();
 sg13g2_fill_8 FILLER_0_67_24 ();
 sg13g2_fill_8 FILLER_0_67_32 ();
 sg13g2_fill_8 FILLER_0_67_40 ();
 sg13g2_fill_8 FILLER_0_67_48 ();
 sg13g2_fill_8 FILLER_0_67_56 ();
 sg13g2_fill_8 FILLER_0_67_64 ();
 sg13g2_fill_8 FILLER_0_67_72 ();
 sg13g2_fill_8 FILLER_0_67_80 ();
 sg13g2_fill_8 FILLER_0_67_88 ();
 sg13g2_fill_8 FILLER_0_67_96 ();
 sg13g2_fill_8 FILLER_0_67_104 ();
 sg13g2_fill_8 FILLER_0_67_112 ();
 sg13g2_fill_8 FILLER_0_67_120 ();
 sg13g2_fill_8 FILLER_0_67_128 ();
 sg13g2_fill_8 FILLER_0_67_136 ();
 sg13g2_fill_8 FILLER_0_67_144 ();
 sg13g2_fill_8 FILLER_0_67_152 ();
 sg13g2_fill_8 FILLER_0_67_160 ();
 sg13g2_fill_8 FILLER_0_67_168 ();
 sg13g2_fill_8 FILLER_0_67_176 ();
 sg13g2_fill_8 FILLER_0_67_184 ();
 sg13g2_fill_8 FILLER_0_67_192 ();
 sg13g2_fill_8 FILLER_0_67_200 ();
 sg13g2_fill_8 FILLER_0_67_208 ();
 sg13g2_fill_8 FILLER_0_67_216 ();
 sg13g2_fill_8 FILLER_0_67_224 ();
 sg13g2_fill_8 FILLER_0_67_232 ();
 sg13g2_fill_8 FILLER_0_67_240 ();
 sg13g2_fill_8 FILLER_0_67_248 ();
 sg13g2_fill_8 FILLER_0_67_256 ();
 sg13g2_fill_8 FILLER_0_67_264 ();
 sg13g2_fill_4 FILLER_0_67_272 ();
 sg13g2_fill_2 FILLER_0_67_276 ();
 sg13g2_fill_1 FILLER_0_67_278 ();
 sg13g2_fill_4 FILLER_0_67_284 ();
 sg13g2_fill_1 FILLER_0_67_288 ();
 sg13g2_fill_2 FILLER_0_67_293 ();
 sg13g2_fill_8 FILLER_0_67_321 ();
 sg13g2_fill_8 FILLER_0_67_329 ();
 sg13g2_fill_8 FILLER_0_67_337 ();
 sg13g2_fill_8 FILLER_0_67_345 ();
 sg13g2_fill_8 FILLER_0_67_353 ();
 sg13g2_fill_2 FILLER_0_67_361 ();
 sg13g2_fill_2 FILLER_0_67_368 ();
 sg13g2_fill_4 FILLER_0_67_375 ();
 sg13g2_fill_1 FILLER_0_67_379 ();
 sg13g2_fill_4 FILLER_0_67_406 ();
 sg13g2_fill_8 FILLER_0_67_416 ();
 sg13g2_fill_4 FILLER_0_67_424 ();
 sg13g2_fill_1 FILLER_0_67_428 ();
 sg13g2_fill_2 FILLER_0_67_434 ();
 sg13g2_fill_4 FILLER_0_67_462 ();
 sg13g2_fill_8 FILLER_0_67_471 ();
 sg13g2_fill_2 FILLER_0_67_484 ();
 sg13g2_fill_2 FILLER_0_67_490 ();
 sg13g2_fill_2 FILLER_0_67_502 ();
 sg13g2_fill_2 FILLER_0_67_530 ();
 sg13g2_fill_2 FILLER_0_67_537 ();
 sg13g2_fill_8 FILLER_0_67_543 ();
 sg13g2_fill_8 FILLER_0_67_551 ();
 sg13g2_fill_8 FILLER_0_67_559 ();
 sg13g2_fill_8 FILLER_0_67_567 ();
 sg13g2_fill_8 FILLER_0_67_575 ();
 sg13g2_fill_8 FILLER_0_67_583 ();
 sg13g2_fill_8 FILLER_0_67_591 ();
 sg13g2_fill_2 FILLER_0_67_599 ();
 sg13g2_fill_1 FILLER_0_67_601 ();
 sg13g2_fill_4 FILLER_0_67_628 ();
 sg13g2_fill_2 FILLER_0_67_632 ();
 sg13g2_fill_1 FILLER_0_67_634 ();
 sg13g2_fill_8 FILLER_0_67_640 ();
 sg13g2_fill_8 FILLER_0_67_652 ();
 sg13g2_fill_4 FILLER_0_67_660 ();
 sg13g2_fill_2 FILLER_0_67_664 ();
 sg13g2_fill_1 FILLER_0_67_666 ();
 sg13g2_fill_4 FILLER_0_67_672 ();
 sg13g2_fill_8 FILLER_0_67_681 ();
 sg13g2_fill_2 FILLER_0_67_689 ();
 sg13g2_fill_1 FILLER_0_67_691 ();
 sg13g2_fill_4 FILLER_0_67_718 ();
 sg13g2_fill_2 FILLER_0_67_726 ();
 sg13g2_fill_1 FILLER_0_67_728 ();
 sg13g2_fill_4 FILLER_0_67_739 ();
 sg13g2_fill_1 FILLER_0_67_743 ();
 sg13g2_fill_2 FILLER_0_67_749 ();
 sg13g2_fill_1 FILLER_0_67_751 ();
 sg13g2_fill_8 FILLER_0_67_778 ();
 sg13g2_fill_8 FILLER_0_67_786 ();
 sg13g2_fill_8 FILLER_0_67_794 ();
 sg13g2_fill_8 FILLER_0_67_802 ();
 sg13g2_fill_8 FILLER_0_67_810 ();
 sg13g2_fill_8 FILLER_0_67_818 ();
 sg13g2_fill_8 FILLER_0_67_826 ();
 sg13g2_fill_4 FILLER_0_67_834 ();
 sg13g2_fill_2 FILLER_0_67_838 ();
 sg13g2_fill_2 FILLER_0_67_845 ();
 sg13g2_fill_8 FILLER_0_67_853 ();
 sg13g2_fill_8 FILLER_0_67_861 ();
 sg13g2_fill_8 FILLER_0_67_869 ();
 sg13g2_fill_8 FILLER_0_67_877 ();
 sg13g2_fill_4 FILLER_0_67_885 ();
 sg13g2_fill_2 FILLER_0_67_894 ();
 sg13g2_fill_8 FILLER_0_67_903 ();
 sg13g2_fill_8 FILLER_0_67_911 ();
 sg13g2_fill_8 FILLER_0_67_919 ();
 sg13g2_fill_1 FILLER_0_67_927 ();
 sg13g2_fill_2 FILLER_0_67_932 ();
 sg13g2_fill_8 FILLER_0_67_944 ();
 sg13g2_fill_8 FILLER_0_67_952 ();
 sg13g2_fill_1 FILLER_0_67_960 ();
 sg13g2_fill_4 FILLER_0_67_966 ();
 sg13g2_fill_1 FILLER_0_67_970 ();
 sg13g2_fill_2 FILLER_0_67_975 ();
 sg13g2_fill_8 FILLER_0_67_981 ();
 sg13g2_fill_8 FILLER_0_67_994 ();
 sg13g2_fill_4 FILLER_0_67_1002 ();
 sg13g2_fill_1 FILLER_0_67_1006 ();
 sg13g2_fill_8 FILLER_0_67_1012 ();
 sg13g2_fill_4 FILLER_0_67_1020 ();
 sg13g2_fill_2 FILLER_0_67_1024 ();
 sg13g2_fill_1 FILLER_0_67_1026 ();
 sg13g2_fill_4 FILLER_0_67_1033 ();
 sg13g2_fill_1 FILLER_0_67_1037 ();
 sg13g2_fill_2 FILLER_0_67_1042 ();
 sg13g2_fill_1 FILLER_0_67_1044 ();
 sg13g2_fill_4 FILLER_0_67_1050 ();
 sg13g2_fill_2 FILLER_0_67_1054 ();
 sg13g2_fill_8 FILLER_0_67_1062 ();
 sg13g2_fill_8 FILLER_0_67_1070 ();
 sg13g2_fill_8 FILLER_0_67_1078 ();
 sg13g2_fill_8 FILLER_0_67_1086 ();
 sg13g2_fill_8 FILLER_0_67_1094 ();
 sg13g2_fill_2 FILLER_0_67_1102 ();
 sg13g2_fill_1 FILLER_0_67_1104 ();
 sg13g2_fill_8 FILLER_0_67_1113 ();
 sg13g2_fill_1 FILLER_0_67_1121 ();
 sg13g2_fill_4 FILLER_0_67_1129 ();
 sg13g2_fill_1 FILLER_0_67_1133 ();
 sg13g2_fill_4 FILLER_0_67_1139 ();
 sg13g2_fill_1 FILLER_0_67_1143 ();
 sg13g2_fill_2 FILLER_0_67_1149 ();
 sg13g2_fill_1 FILLER_0_67_1151 ();
 sg13g2_fill_2 FILLER_0_67_1157 ();
 sg13g2_fill_8 FILLER_0_67_1164 ();
 sg13g2_fill_1 FILLER_0_67_1172 ();
 sg13g2_fill_8 FILLER_0_67_1181 ();
 sg13g2_fill_8 FILLER_0_67_1189 ();
 sg13g2_fill_8 FILLER_0_67_1197 ();
 sg13g2_fill_8 FILLER_0_67_1210 ();
 sg13g2_fill_4 FILLER_0_67_1218 ();
 sg13g2_fill_2 FILLER_0_67_1222 ();
 sg13g2_fill_1 FILLER_0_67_1224 ();
 sg13g2_fill_2 FILLER_0_67_1229 ();
 sg13g2_fill_8 FILLER_0_67_1236 ();
 sg13g2_fill_8 FILLER_0_67_1244 ();
 sg13g2_fill_8 FILLER_0_67_1252 ();
 sg13g2_fill_8 FILLER_0_67_1260 ();
 sg13g2_fill_4 FILLER_0_67_1268 ();
 sg13g2_fill_1 FILLER_0_67_1272 ();
 sg13g2_fill_2 FILLER_0_67_1278 ();
 sg13g2_fill_8 FILLER_0_67_1285 ();
 sg13g2_fill_4 FILLER_0_67_1293 ();
 sg13g2_fill_8 FILLER_0_68_0 ();
 sg13g2_fill_8 FILLER_0_68_8 ();
 sg13g2_fill_8 FILLER_0_68_16 ();
 sg13g2_fill_8 FILLER_0_68_24 ();
 sg13g2_fill_8 FILLER_0_68_32 ();
 sg13g2_fill_8 FILLER_0_68_40 ();
 sg13g2_fill_8 FILLER_0_68_48 ();
 sg13g2_fill_8 FILLER_0_68_56 ();
 sg13g2_fill_8 FILLER_0_68_64 ();
 sg13g2_fill_8 FILLER_0_68_72 ();
 sg13g2_fill_8 FILLER_0_68_80 ();
 sg13g2_fill_8 FILLER_0_68_88 ();
 sg13g2_fill_8 FILLER_0_68_96 ();
 sg13g2_fill_8 FILLER_0_68_104 ();
 sg13g2_fill_8 FILLER_0_68_112 ();
 sg13g2_fill_8 FILLER_0_68_120 ();
 sg13g2_fill_8 FILLER_0_68_128 ();
 sg13g2_fill_8 FILLER_0_68_136 ();
 sg13g2_fill_8 FILLER_0_68_144 ();
 sg13g2_fill_8 FILLER_0_68_152 ();
 sg13g2_fill_8 FILLER_0_68_160 ();
 sg13g2_fill_8 FILLER_0_68_168 ();
 sg13g2_fill_8 FILLER_0_68_176 ();
 sg13g2_fill_8 FILLER_0_68_184 ();
 sg13g2_fill_8 FILLER_0_68_192 ();
 sg13g2_fill_4 FILLER_0_68_200 ();
 sg13g2_fill_2 FILLER_0_68_204 ();
 sg13g2_fill_1 FILLER_0_68_206 ();
 sg13g2_fill_2 FILLER_0_68_233 ();
 sg13g2_fill_8 FILLER_0_68_240 ();
 sg13g2_fill_2 FILLER_0_68_254 ();
 sg13g2_fill_8 FILLER_0_68_261 ();
 sg13g2_fill_8 FILLER_0_68_269 ();
 sg13g2_fill_8 FILLER_0_68_277 ();
 sg13g2_fill_8 FILLER_0_68_285 ();
 sg13g2_fill_8 FILLER_0_68_293 ();
 sg13g2_fill_8 FILLER_0_68_301 ();
 sg13g2_fill_4 FILLER_0_68_309 ();
 sg13g2_fill_2 FILLER_0_68_313 ();
 sg13g2_fill_1 FILLER_0_68_315 ();
 sg13g2_fill_8 FILLER_0_68_321 ();
 sg13g2_fill_8 FILLER_0_68_329 ();
 sg13g2_fill_8 FILLER_0_68_337 ();
 sg13g2_fill_8 FILLER_0_68_345 ();
 sg13g2_fill_4 FILLER_0_68_353 ();
 sg13g2_fill_4 FILLER_0_68_362 ();
 sg13g2_fill_2 FILLER_0_68_366 ();
 sg13g2_fill_8 FILLER_0_68_376 ();
 sg13g2_fill_8 FILLER_0_68_384 ();
 sg13g2_fill_2 FILLER_0_68_392 ();
 sg13g2_fill_2 FILLER_0_68_399 ();
 sg13g2_fill_4 FILLER_0_68_405 ();
 sg13g2_fill_1 FILLER_0_68_409 ();
 sg13g2_fill_8 FILLER_0_68_415 ();
 sg13g2_fill_8 FILLER_0_68_423 ();
 sg13g2_fill_1 FILLER_0_68_431 ();
 sg13g2_fill_8 FILLER_0_68_437 ();
 sg13g2_fill_4 FILLER_0_68_445 ();
 sg13g2_fill_2 FILLER_0_68_449 ();
 sg13g2_fill_1 FILLER_0_68_451 ();
 sg13g2_fill_2 FILLER_0_68_456 ();
 sg13g2_fill_2 FILLER_0_68_468 ();
 sg13g2_fill_8 FILLER_0_68_475 ();
 sg13g2_fill_8 FILLER_0_68_483 ();
 sg13g2_fill_8 FILLER_0_68_491 ();
 sg13g2_fill_8 FILLER_0_68_499 ();
 sg13g2_fill_4 FILLER_0_68_507 ();
 sg13g2_fill_8 FILLER_0_68_516 ();
 sg13g2_fill_8 FILLER_0_68_524 ();
 sg13g2_fill_8 FILLER_0_68_532 ();
 sg13g2_fill_8 FILLER_0_68_540 ();
 sg13g2_fill_1 FILLER_0_68_548 ();
 sg13g2_fill_2 FILLER_0_68_553 ();
 sg13g2_fill_2 FILLER_0_68_581 ();
 sg13g2_fill_8 FILLER_0_68_593 ();
 sg13g2_fill_8 FILLER_0_68_601 ();
 sg13g2_fill_8 FILLER_0_68_609 ();
 sg13g2_fill_8 FILLER_0_68_617 ();
 sg13g2_fill_8 FILLER_0_68_625 ();
 sg13g2_fill_8 FILLER_0_68_633 ();
 sg13g2_fill_8 FILLER_0_68_641 ();
 sg13g2_fill_4 FILLER_0_68_649 ();
 sg13g2_fill_2 FILLER_0_68_657 ();
 sg13g2_fill_2 FILLER_0_68_664 ();
 sg13g2_fill_4 FILLER_0_68_670 ();
 sg13g2_fill_2 FILLER_0_68_674 ();
 sg13g2_fill_8 FILLER_0_68_682 ();
 sg13g2_fill_1 FILLER_0_68_690 ();
 sg13g2_fill_4 FILLER_0_68_701 ();
 sg13g2_fill_1 FILLER_0_68_705 ();
 sg13g2_fill_8 FILLER_0_68_732 ();
 sg13g2_fill_1 FILLER_0_68_740 ();
 sg13g2_fill_2 FILLER_0_68_747 ();
 sg13g2_fill_2 FILLER_0_68_759 ();
 sg13g2_fill_2 FILLER_0_68_766 ();
 sg13g2_fill_2 FILLER_0_68_774 ();
 sg13g2_fill_8 FILLER_0_68_781 ();
 sg13g2_fill_2 FILLER_0_68_789 ();
 sg13g2_fill_8 FILLER_0_68_801 ();
 sg13g2_fill_4 FILLER_0_68_809 ();
 sg13g2_fill_8 FILLER_0_68_823 ();
 sg13g2_fill_8 FILLER_0_68_837 ();
 sg13g2_fill_8 FILLER_0_68_845 ();
 sg13g2_fill_8 FILLER_0_68_853 ();
 sg13g2_fill_8 FILLER_0_68_861 ();
 sg13g2_fill_8 FILLER_0_68_869 ();
 sg13g2_fill_1 FILLER_0_68_877 ();
 sg13g2_fill_2 FILLER_0_68_882 ();
 sg13g2_fill_2 FILLER_0_68_889 ();
 sg13g2_fill_8 FILLER_0_68_901 ();
 sg13g2_fill_4 FILLER_0_68_909 ();
 sg13g2_fill_2 FILLER_0_68_913 ();
 sg13g2_fill_2 FILLER_0_68_925 ();
 sg13g2_fill_4 FILLER_0_68_933 ();
 sg13g2_fill_4 FILLER_0_68_943 ();
 sg13g2_fill_1 FILLER_0_68_947 ();
 sg13g2_fill_8 FILLER_0_68_954 ();
 sg13g2_fill_4 FILLER_0_68_967 ();
 sg13g2_fill_4 FILLER_0_68_976 ();
 sg13g2_fill_2 FILLER_0_68_984 ();
 sg13g2_fill_8 FILLER_0_68_992 ();
 sg13g2_fill_1 FILLER_0_68_1000 ();
 sg13g2_fill_4 FILLER_0_68_1007 ();
 sg13g2_fill_2 FILLER_0_68_1011 ();
 sg13g2_fill_1 FILLER_0_68_1013 ();
 sg13g2_fill_8 FILLER_0_68_1019 ();
 sg13g2_fill_1 FILLER_0_68_1027 ();
 sg13g2_fill_2 FILLER_0_68_1033 ();
 sg13g2_fill_2 FILLER_0_68_1041 ();
 sg13g2_fill_4 FILLER_0_68_1048 ();
 sg13g2_fill_2 FILLER_0_68_1052 ();
 sg13g2_fill_8 FILLER_0_68_1061 ();
 sg13g2_fill_8 FILLER_0_68_1069 ();
 sg13g2_fill_8 FILLER_0_68_1077 ();
 sg13g2_fill_2 FILLER_0_68_1085 ();
 sg13g2_fill_1 FILLER_0_68_1087 ();
 sg13g2_fill_8 FILLER_0_68_1092 ();
 sg13g2_fill_4 FILLER_0_68_1100 ();
 sg13g2_fill_2 FILLER_0_68_1104 ();
 sg13g2_fill_1 FILLER_0_68_1106 ();
 sg13g2_fill_4 FILLER_0_68_1114 ();
 sg13g2_fill_2 FILLER_0_68_1123 ();
 sg13g2_fill_8 FILLER_0_68_1130 ();
 sg13g2_fill_8 FILLER_0_68_1138 ();
 sg13g2_fill_8 FILLER_0_68_1146 ();
 sg13g2_fill_8 FILLER_0_68_1154 ();
 sg13g2_fill_1 FILLER_0_68_1162 ();
 sg13g2_fill_8 FILLER_0_68_1171 ();
 sg13g2_fill_8 FILLER_0_68_1179 ();
 sg13g2_fill_8 FILLER_0_68_1187 ();
 sg13g2_fill_4 FILLER_0_68_1195 ();
 sg13g2_fill_2 FILLER_0_68_1199 ();
 sg13g2_fill_1 FILLER_0_68_1201 ();
 sg13g2_fill_2 FILLER_0_68_1207 ();
 sg13g2_fill_2 FILLER_0_68_1214 ();
 sg13g2_fill_1 FILLER_0_68_1216 ();
 sg13g2_fill_2 FILLER_0_68_1222 ();
 sg13g2_fill_2 FILLER_0_68_1228 ();
 sg13g2_fill_8 FILLER_0_68_1235 ();
 sg13g2_fill_8 FILLER_0_68_1243 ();
 sg13g2_fill_2 FILLER_0_68_1261 ();
 sg13g2_fill_8 FILLER_0_68_1289 ();
 sg13g2_fill_8 FILLER_0_69_0 ();
 sg13g2_fill_8 FILLER_0_69_8 ();
 sg13g2_fill_8 FILLER_0_69_16 ();
 sg13g2_fill_8 FILLER_0_69_24 ();
 sg13g2_fill_8 FILLER_0_69_32 ();
 sg13g2_fill_8 FILLER_0_69_40 ();
 sg13g2_fill_8 FILLER_0_69_48 ();
 sg13g2_fill_8 FILLER_0_69_56 ();
 sg13g2_fill_8 FILLER_0_69_64 ();
 sg13g2_fill_8 FILLER_0_69_72 ();
 sg13g2_fill_8 FILLER_0_69_80 ();
 sg13g2_fill_8 FILLER_0_69_88 ();
 sg13g2_fill_8 FILLER_0_69_96 ();
 sg13g2_fill_8 FILLER_0_69_104 ();
 sg13g2_fill_8 FILLER_0_69_112 ();
 sg13g2_fill_8 FILLER_0_69_120 ();
 sg13g2_fill_8 FILLER_0_69_128 ();
 sg13g2_fill_8 FILLER_0_69_136 ();
 sg13g2_fill_8 FILLER_0_69_144 ();
 sg13g2_fill_8 FILLER_0_69_152 ();
 sg13g2_fill_8 FILLER_0_69_160 ();
 sg13g2_fill_8 FILLER_0_69_168 ();
 sg13g2_fill_8 FILLER_0_69_176 ();
 sg13g2_fill_8 FILLER_0_69_184 ();
 sg13g2_fill_8 FILLER_0_69_192 ();
 sg13g2_fill_8 FILLER_0_69_200 ();
 sg13g2_fill_4 FILLER_0_69_213 ();
 sg13g2_fill_2 FILLER_0_69_217 ();
 sg13g2_fill_8 FILLER_0_69_245 ();
 sg13g2_fill_8 FILLER_0_69_253 ();
 sg13g2_fill_8 FILLER_0_69_261 ();
 sg13g2_fill_1 FILLER_0_69_269 ();
 sg13g2_fill_4 FILLER_0_69_296 ();
 sg13g2_fill_2 FILLER_0_69_300 ();
 sg13g2_fill_1 FILLER_0_69_302 ();
 sg13g2_fill_8 FILLER_0_69_307 ();
 sg13g2_fill_8 FILLER_0_69_315 ();
 sg13g2_fill_8 FILLER_0_69_323 ();
 sg13g2_fill_8 FILLER_0_69_331 ();
 sg13g2_fill_2 FILLER_0_69_339 ();
 sg13g2_fill_1 FILLER_0_69_341 ();
 sg13g2_fill_2 FILLER_0_69_347 ();
 sg13g2_fill_8 FILLER_0_69_357 ();
 sg13g2_fill_8 FILLER_0_69_365 ();
 sg13g2_fill_8 FILLER_0_69_373 ();
 sg13g2_fill_8 FILLER_0_69_381 ();
 sg13g2_fill_8 FILLER_0_69_389 ();
 sg13g2_fill_8 FILLER_0_69_397 ();
 sg13g2_fill_8 FILLER_0_69_405 ();
 sg13g2_fill_8 FILLER_0_69_413 ();
 sg13g2_fill_8 FILLER_0_69_421 ();
 sg13g2_fill_8 FILLER_0_69_429 ();
 sg13g2_fill_8 FILLER_0_69_437 ();
 sg13g2_fill_8 FILLER_0_69_445 ();
 sg13g2_fill_8 FILLER_0_69_453 ();
 sg13g2_fill_8 FILLER_0_69_461 ();
 sg13g2_fill_4 FILLER_0_69_469 ();
 sg13g2_fill_2 FILLER_0_69_473 ();
 sg13g2_fill_1 FILLER_0_69_475 ();
 sg13g2_fill_8 FILLER_0_69_481 ();
 sg13g2_fill_8 FILLER_0_69_489 ();
 sg13g2_fill_2 FILLER_0_69_497 ();
 sg13g2_fill_4 FILLER_0_69_504 ();
 sg13g2_fill_2 FILLER_0_69_508 ();
 sg13g2_fill_2 FILLER_0_69_515 ();
 sg13g2_fill_2 FILLER_0_69_522 ();
 sg13g2_fill_1 FILLER_0_69_524 ();
 sg13g2_fill_8 FILLER_0_69_529 ();
 sg13g2_fill_4 FILLER_0_69_537 ();
 sg13g2_fill_2 FILLER_0_69_541 ();
 sg13g2_fill_2 FILLER_0_69_548 ();
 sg13g2_fill_2 FILLER_0_69_555 ();
 sg13g2_fill_2 FILLER_0_69_583 ();
 sg13g2_fill_4 FILLER_0_69_590 ();
 sg13g2_fill_1 FILLER_0_69_594 ();
 sg13g2_fill_2 FILLER_0_69_600 ();
 sg13g2_fill_8 FILLER_0_69_607 ();
 sg13g2_fill_4 FILLER_0_69_615 ();
 sg13g2_fill_2 FILLER_0_69_624 ();
 sg13g2_fill_1 FILLER_0_69_626 ();
 sg13g2_fill_4 FILLER_0_69_631 ();
 sg13g2_fill_2 FILLER_0_69_635 ();
 sg13g2_fill_8 FILLER_0_69_643 ();
 sg13g2_fill_4 FILLER_0_69_651 ();
 sg13g2_fill_2 FILLER_0_69_655 ();
 sg13g2_fill_8 FILLER_0_69_683 ();
 sg13g2_fill_8 FILLER_0_69_691 ();
 sg13g2_fill_4 FILLER_0_69_709 ();
 sg13g2_fill_2 FILLER_0_69_713 ();
 sg13g2_fill_8 FILLER_0_69_725 ();
 sg13g2_fill_8 FILLER_0_69_738 ();
 sg13g2_fill_8 FILLER_0_69_746 ();
 sg13g2_fill_2 FILLER_0_69_754 ();
 sg13g2_fill_8 FILLER_0_69_761 ();
 sg13g2_fill_1 FILLER_0_69_769 ();
 sg13g2_fill_2 FILLER_0_69_775 ();
 sg13g2_fill_2 FILLER_0_69_783 ();
 sg13g2_fill_4 FILLER_0_69_811 ();
 sg13g2_fill_1 FILLER_0_69_815 ();
 sg13g2_fill_8 FILLER_0_69_842 ();
 sg13g2_fill_8 FILLER_0_69_850 ();
 sg13g2_fill_4 FILLER_0_69_858 ();
 sg13g2_fill_1 FILLER_0_69_862 ();
 sg13g2_fill_2 FILLER_0_69_871 ();
 sg13g2_fill_2 FILLER_0_69_877 ();
 sg13g2_fill_4 FILLER_0_69_884 ();
 sg13g2_fill_2 FILLER_0_69_893 ();
 sg13g2_fill_8 FILLER_0_69_916 ();
 sg13g2_fill_8 FILLER_0_69_924 ();
 sg13g2_fill_2 FILLER_0_69_932 ();
 sg13g2_fill_2 FILLER_0_69_939 ();
 sg13g2_fill_2 FILLER_0_69_945 ();
 sg13g2_fill_2 FILLER_0_69_952 ();
 sg13g2_fill_8 FILLER_0_69_958 ();
 sg13g2_fill_2 FILLER_0_69_966 ();
 sg13g2_fill_1 FILLER_0_69_968 ();
 sg13g2_fill_2 FILLER_0_69_974 ();
 sg13g2_fill_2 FILLER_0_69_980 ();
 sg13g2_fill_2 FILLER_0_69_986 ();
 sg13g2_fill_2 FILLER_0_69_994 ();
 sg13g2_fill_4 FILLER_0_69_1001 ();
 sg13g2_fill_2 FILLER_0_69_1005 ();
 sg13g2_fill_2 FILLER_0_69_1012 ();
 sg13g2_fill_2 FILLER_0_69_1020 ();
 sg13g2_fill_4 FILLER_0_69_1027 ();
 sg13g2_fill_2 FILLER_0_69_1031 ();
 sg13g2_fill_1 FILLER_0_69_1033 ();
 sg13g2_fill_4 FILLER_0_69_1039 ();
 sg13g2_fill_2 FILLER_0_69_1043 ();
 sg13g2_fill_1 FILLER_0_69_1045 ();
 sg13g2_fill_2 FILLER_0_69_1050 ();
 sg13g2_fill_2 FILLER_0_69_1056 ();
 sg13g2_fill_1 FILLER_0_69_1058 ();
 sg13g2_fill_8 FILLER_0_69_1065 ();
 sg13g2_fill_8 FILLER_0_69_1073 ();
 sg13g2_fill_8 FILLER_0_69_1081 ();
 sg13g2_fill_8 FILLER_0_69_1089 ();
 sg13g2_fill_1 FILLER_0_69_1097 ();
 sg13g2_fill_2 FILLER_0_69_1103 ();
 sg13g2_fill_2 FILLER_0_69_1110 ();
 sg13g2_fill_8 FILLER_0_69_1117 ();
 sg13g2_fill_8 FILLER_0_69_1125 ();
 sg13g2_fill_4 FILLER_0_69_1133 ();
 sg13g2_fill_1 FILLER_0_69_1137 ();
 sg13g2_fill_8 FILLER_0_69_1142 ();
 sg13g2_fill_2 FILLER_0_69_1150 ();
 sg13g2_fill_2 FILLER_0_69_1156 ();
 sg13g2_fill_1 FILLER_0_69_1158 ();
 sg13g2_fill_2 FILLER_0_69_1164 ();
 sg13g2_fill_8 FILLER_0_69_1171 ();
 sg13g2_fill_1 FILLER_0_69_1179 ();
 sg13g2_fill_8 FILLER_0_69_1188 ();
 sg13g2_fill_8 FILLER_0_69_1196 ();
 sg13g2_fill_4 FILLER_0_69_1204 ();
 sg13g2_fill_1 FILLER_0_69_1208 ();
 sg13g2_fill_2 FILLER_0_69_1213 ();
 sg13g2_fill_1 FILLER_0_69_1215 ();
 sg13g2_fill_4 FILLER_0_69_1224 ();
 sg13g2_fill_4 FILLER_0_69_1233 ();
 sg13g2_fill_1 FILLER_0_69_1237 ();
 sg13g2_fill_4 FILLER_0_69_1246 ();
 sg13g2_fill_2 FILLER_0_69_1250 ();
 sg13g2_fill_1 FILLER_0_69_1252 ();
 sg13g2_fill_2 FILLER_0_69_1263 ();
 sg13g2_fill_8 FILLER_0_69_1270 ();
 sg13g2_fill_1 FILLER_0_69_1278 ();
 sg13g2_fill_8 FILLER_0_69_1287 ();
 sg13g2_fill_2 FILLER_0_69_1295 ();
 sg13g2_fill_8 FILLER_0_70_0 ();
 sg13g2_fill_8 FILLER_0_70_8 ();
 sg13g2_fill_8 FILLER_0_70_16 ();
 sg13g2_fill_8 FILLER_0_70_24 ();
 sg13g2_fill_8 FILLER_0_70_32 ();
 sg13g2_fill_8 FILLER_0_70_40 ();
 sg13g2_fill_8 FILLER_0_70_48 ();
 sg13g2_fill_8 FILLER_0_70_56 ();
 sg13g2_fill_8 FILLER_0_70_64 ();
 sg13g2_fill_8 FILLER_0_70_72 ();
 sg13g2_fill_8 FILLER_0_70_80 ();
 sg13g2_fill_8 FILLER_0_70_88 ();
 sg13g2_fill_8 FILLER_0_70_96 ();
 sg13g2_fill_8 FILLER_0_70_104 ();
 sg13g2_fill_8 FILLER_0_70_112 ();
 sg13g2_fill_8 FILLER_0_70_120 ();
 sg13g2_fill_8 FILLER_0_70_128 ();
 sg13g2_fill_8 FILLER_0_70_136 ();
 sg13g2_fill_8 FILLER_0_70_144 ();
 sg13g2_fill_8 FILLER_0_70_152 ();
 sg13g2_fill_8 FILLER_0_70_160 ();
 sg13g2_fill_8 FILLER_0_70_168 ();
 sg13g2_fill_8 FILLER_0_70_176 ();
 sg13g2_fill_8 FILLER_0_70_184 ();
 sg13g2_fill_8 FILLER_0_70_192 ();
 sg13g2_fill_8 FILLER_0_70_200 ();
 sg13g2_fill_4 FILLER_0_70_208 ();
 sg13g2_fill_2 FILLER_0_70_212 ();
 sg13g2_fill_2 FILLER_0_70_218 ();
 sg13g2_fill_2 FILLER_0_70_225 ();
 sg13g2_fill_4 FILLER_0_70_231 ();
 sg13g2_fill_1 FILLER_0_70_235 ();
 sg13g2_fill_8 FILLER_0_70_257 ();
 sg13g2_fill_8 FILLER_0_70_265 ();
 sg13g2_fill_8 FILLER_0_70_273 ();
 sg13g2_fill_4 FILLER_0_70_281 ();
 sg13g2_fill_1 FILLER_0_70_285 ();
 sg13g2_fill_2 FILLER_0_70_291 ();
 sg13g2_fill_4 FILLER_0_70_298 ();
 sg13g2_fill_1 FILLER_0_70_302 ();
 sg13g2_fill_2 FILLER_0_70_309 ();
 sg13g2_fill_8 FILLER_0_70_316 ();
 sg13g2_fill_2 FILLER_0_70_328 ();
 sg13g2_fill_2 FILLER_0_70_336 ();
 sg13g2_fill_2 FILLER_0_70_345 ();
 sg13g2_fill_2 FILLER_0_70_373 ();
 sg13g2_fill_2 FILLER_0_70_380 ();
 sg13g2_fill_8 FILLER_0_70_386 ();
 sg13g2_fill_8 FILLER_0_70_394 ();
 sg13g2_fill_8 FILLER_0_70_407 ();
 sg13g2_fill_4 FILLER_0_70_419 ();
 sg13g2_fill_2 FILLER_0_70_449 ();
 sg13g2_fill_2 FILLER_0_70_456 ();
 sg13g2_fill_2 FILLER_0_70_463 ();
 sg13g2_fill_8 FILLER_0_70_469 ();
 sg13g2_fill_2 FILLER_0_70_482 ();
 sg13g2_fill_1 FILLER_0_70_484 ();
 sg13g2_fill_4 FILLER_0_70_495 ();
 sg13g2_fill_2 FILLER_0_70_499 ();
 sg13g2_fill_1 FILLER_0_70_501 ();
 sg13g2_fill_4 FILLER_0_70_508 ();
 sg13g2_fill_2 FILLER_0_70_517 ();
 sg13g2_fill_8 FILLER_0_70_524 ();
 sg13g2_fill_2 FILLER_0_70_532 ();
 sg13g2_fill_1 FILLER_0_70_534 ();
 sg13g2_fill_4 FILLER_0_70_545 ();
 sg13g2_fill_1 FILLER_0_70_549 ();
 sg13g2_fill_8 FILLER_0_70_554 ();
 sg13g2_fill_8 FILLER_0_70_562 ();
 sg13g2_fill_8 FILLER_0_70_570 ();
 sg13g2_fill_8 FILLER_0_70_578 ();
 sg13g2_fill_8 FILLER_0_70_586 ();
 sg13g2_fill_4 FILLER_0_70_598 ();
 sg13g2_fill_2 FILLER_0_70_607 ();
 sg13g2_fill_4 FILLER_0_70_635 ();
 sg13g2_fill_2 FILLER_0_70_644 ();
 sg13g2_fill_2 FILLER_0_70_672 ();
 sg13g2_fill_8 FILLER_0_70_679 ();
 sg13g2_fill_8 FILLER_0_70_687 ();
 sg13g2_fill_8 FILLER_0_70_695 ();
 sg13g2_fill_8 FILLER_0_70_703 ();
 sg13g2_fill_1 FILLER_0_70_711 ();
 sg13g2_fill_8 FILLER_0_70_717 ();
 sg13g2_fill_8 FILLER_0_70_725 ();
 sg13g2_fill_2 FILLER_0_70_733 ();
 sg13g2_fill_1 FILLER_0_70_735 ();
 sg13g2_fill_8 FILLER_0_70_742 ();
 sg13g2_fill_8 FILLER_0_70_750 ();
 sg13g2_fill_8 FILLER_0_70_758 ();
 sg13g2_fill_8 FILLER_0_70_766 ();
 sg13g2_fill_8 FILLER_0_70_774 ();
 sg13g2_fill_8 FILLER_0_70_782 ();
 sg13g2_fill_8 FILLER_0_70_790 ();
 sg13g2_fill_8 FILLER_0_70_804 ();
 sg13g2_fill_4 FILLER_0_70_812 ();
 sg13g2_fill_8 FILLER_0_70_826 ();
 sg13g2_fill_8 FILLER_0_70_834 ();
 sg13g2_fill_8 FILLER_0_70_842 ();
 sg13g2_fill_8 FILLER_0_70_850 ();
 sg13g2_fill_4 FILLER_0_70_858 ();
 sg13g2_fill_1 FILLER_0_70_862 ();
 sg13g2_fill_2 FILLER_0_70_871 ();
 sg13g2_fill_2 FILLER_0_70_878 ();
 sg13g2_fill_8 FILLER_0_70_887 ();
 sg13g2_fill_2 FILLER_0_70_895 ();
 sg13g2_fill_8 FILLER_0_70_901 ();
 sg13g2_fill_4 FILLER_0_70_909 ();
 sg13g2_fill_2 FILLER_0_70_913 ();
 sg13g2_fill_2 FILLER_0_70_920 ();
 sg13g2_fill_8 FILLER_0_70_928 ();
 sg13g2_fill_2 FILLER_0_70_936 ();
 sg13g2_fill_1 FILLER_0_70_938 ();
 sg13g2_fill_2 FILLER_0_70_943 ();
 sg13g2_fill_2 FILLER_0_70_950 ();
 sg13g2_fill_8 FILLER_0_70_957 ();
 sg13g2_fill_2 FILLER_0_70_965 ();
 sg13g2_fill_1 FILLER_0_70_967 ();
 sg13g2_fill_4 FILLER_0_70_973 ();
 sg13g2_fill_1 FILLER_0_70_977 ();
 sg13g2_fill_2 FILLER_0_70_988 ();
 sg13g2_fill_4 FILLER_0_70_996 ();
 sg13g2_fill_2 FILLER_0_70_1000 ();
 sg13g2_fill_1 FILLER_0_70_1002 ();
 sg13g2_fill_2 FILLER_0_70_1008 ();
 sg13g2_fill_4 FILLER_0_70_1016 ();
 sg13g2_fill_1 FILLER_0_70_1020 ();
 sg13g2_fill_2 FILLER_0_70_1026 ();
 sg13g2_fill_4 FILLER_0_70_1032 ();
 sg13g2_fill_1 FILLER_0_70_1036 ();
 sg13g2_fill_2 FILLER_0_70_1042 ();
 sg13g2_fill_1 FILLER_0_70_1044 ();
 sg13g2_fill_4 FILLER_0_70_1052 ();
 sg13g2_fill_8 FILLER_0_70_1060 ();
 sg13g2_fill_2 FILLER_0_70_1068 ();
 sg13g2_fill_2 FILLER_0_70_1078 ();
 sg13g2_fill_2 FILLER_0_70_1088 ();
 sg13g2_fill_1 FILLER_0_70_1090 ();
 sg13g2_fill_4 FILLER_0_70_1096 ();
 sg13g2_fill_2 FILLER_0_70_1100 ();
 sg13g2_fill_1 FILLER_0_70_1102 ();
 sg13g2_fill_4 FILLER_0_70_1106 ();
 sg13g2_fill_2 FILLER_0_70_1110 ();
 sg13g2_fill_8 FILLER_0_70_1117 ();
 sg13g2_fill_8 FILLER_0_70_1125 ();
 sg13g2_fill_4 FILLER_0_70_1133 ();
 sg13g2_fill_2 FILLER_0_70_1137 ();
 sg13g2_fill_1 FILLER_0_70_1139 ();
 sg13g2_fill_8 FILLER_0_70_1145 ();
 sg13g2_fill_4 FILLER_0_70_1153 ();
 sg13g2_fill_4 FILLER_0_70_1165 ();
 sg13g2_fill_4 FILLER_0_70_1173 ();
 sg13g2_fill_4 FILLER_0_70_1181 ();
 sg13g2_fill_8 FILLER_0_70_1190 ();
 sg13g2_fill_8 FILLER_0_70_1198 ();
 sg13g2_fill_8 FILLER_0_70_1206 ();
 sg13g2_fill_4 FILLER_0_70_1214 ();
 sg13g2_fill_2 FILLER_0_70_1218 ();
 sg13g2_fill_1 FILLER_0_70_1220 ();
 sg13g2_fill_2 FILLER_0_70_1228 ();
 sg13g2_fill_4 FILLER_0_70_1235 ();
 sg13g2_fill_2 FILLER_0_70_1244 ();
 sg13g2_fill_1 FILLER_0_70_1246 ();
 sg13g2_fill_8 FILLER_0_70_1252 ();
 sg13g2_fill_1 FILLER_0_70_1260 ();
 sg13g2_fill_2 FILLER_0_70_1269 ();
 sg13g2_fill_4 FILLER_0_70_1275 ();
 sg13g2_fill_2 FILLER_0_70_1279 ();
 sg13g2_fill_2 FILLER_0_70_1285 ();
 sg13g2_fill_4 FILLER_0_70_1292 ();
 sg13g2_fill_1 FILLER_0_70_1296 ();
 sg13g2_fill_8 FILLER_0_71_0 ();
 sg13g2_fill_8 FILLER_0_71_8 ();
 sg13g2_fill_8 FILLER_0_71_16 ();
 sg13g2_fill_8 FILLER_0_71_24 ();
 sg13g2_fill_8 FILLER_0_71_32 ();
 sg13g2_fill_8 FILLER_0_71_40 ();
 sg13g2_fill_8 FILLER_0_71_48 ();
 sg13g2_fill_8 FILLER_0_71_56 ();
 sg13g2_fill_8 FILLER_0_71_64 ();
 sg13g2_fill_8 FILLER_0_71_72 ();
 sg13g2_fill_8 FILLER_0_71_80 ();
 sg13g2_fill_8 FILLER_0_71_88 ();
 sg13g2_fill_8 FILLER_0_71_96 ();
 sg13g2_fill_8 FILLER_0_71_104 ();
 sg13g2_fill_8 FILLER_0_71_112 ();
 sg13g2_fill_8 FILLER_0_71_120 ();
 sg13g2_fill_8 FILLER_0_71_128 ();
 sg13g2_fill_8 FILLER_0_71_136 ();
 sg13g2_fill_8 FILLER_0_71_144 ();
 sg13g2_fill_8 FILLER_0_71_152 ();
 sg13g2_fill_8 FILLER_0_71_160 ();
 sg13g2_fill_8 FILLER_0_71_168 ();
 sg13g2_fill_8 FILLER_0_71_176 ();
 sg13g2_fill_8 FILLER_0_71_184 ();
 sg13g2_fill_8 FILLER_0_71_192 ();
 sg13g2_fill_8 FILLER_0_71_200 ();
 sg13g2_fill_8 FILLER_0_71_208 ();
 sg13g2_fill_8 FILLER_0_71_216 ();
 sg13g2_fill_2 FILLER_0_71_224 ();
 sg13g2_fill_8 FILLER_0_71_230 ();
 sg13g2_fill_4 FILLER_0_71_238 ();
 sg13g2_fill_2 FILLER_0_71_242 ();
 sg13g2_fill_4 FILLER_0_71_249 ();
 sg13g2_fill_1 FILLER_0_71_253 ();
 sg13g2_fill_8 FILLER_0_71_258 ();
 sg13g2_fill_8 FILLER_0_71_266 ();
 sg13g2_fill_4 FILLER_0_71_274 ();
 sg13g2_fill_2 FILLER_0_71_304 ();
 sg13g2_fill_2 FILLER_0_71_312 ();
 sg13g2_fill_4 FILLER_0_71_340 ();
 sg13g2_fill_4 FILLER_0_71_348 ();
 sg13g2_fill_2 FILLER_0_71_352 ();
 sg13g2_fill_1 FILLER_0_71_354 ();
 sg13g2_fill_2 FILLER_0_71_360 ();
 sg13g2_fill_1 FILLER_0_71_362 ();
 sg13g2_fill_4 FILLER_0_71_389 ();
 sg13g2_fill_2 FILLER_0_71_393 ();
 sg13g2_fill_1 FILLER_0_71_395 ();
 sg13g2_fill_2 FILLER_0_71_422 ();
 sg13g2_fill_2 FILLER_0_71_429 ();
 sg13g2_fill_1 FILLER_0_71_431 ();
 sg13g2_fill_2 FILLER_0_71_437 ();
 sg13g2_fill_1 FILLER_0_71_439 ();
 sg13g2_fill_2 FILLER_0_71_466 ();
 sg13g2_fill_1 FILLER_0_71_468 ();
 sg13g2_fill_2 FILLER_0_71_495 ();
 sg13g2_fill_1 FILLER_0_71_497 ();
 sg13g2_fill_4 FILLER_0_71_502 ();
 sg13g2_fill_2 FILLER_0_71_506 ();
 sg13g2_fill_1 FILLER_0_71_508 ();
 sg13g2_fill_8 FILLER_0_71_535 ();
 sg13g2_fill_1 FILLER_0_71_543 ();
 sg13g2_fill_8 FILLER_0_71_549 ();
 sg13g2_fill_8 FILLER_0_71_557 ();
 sg13g2_fill_8 FILLER_0_71_565 ();
 sg13g2_fill_8 FILLER_0_71_573 ();
 sg13g2_fill_8 FILLER_0_71_581 ();
 sg13g2_fill_8 FILLER_0_71_589 ();
 sg13g2_fill_4 FILLER_0_71_597 ();
 sg13g2_fill_2 FILLER_0_71_601 ();
 sg13g2_fill_8 FILLER_0_71_608 ();
 sg13g2_fill_8 FILLER_0_71_616 ();
 sg13g2_fill_8 FILLER_0_71_624 ();
 sg13g2_fill_8 FILLER_0_71_632 ();
 sg13g2_fill_8 FILLER_0_71_640 ();
 sg13g2_fill_4 FILLER_0_71_648 ();
 sg13g2_fill_2 FILLER_0_71_652 ();
 sg13g2_fill_1 FILLER_0_71_654 ();
 sg13g2_fill_4 FILLER_0_71_659 ();
 sg13g2_fill_8 FILLER_0_71_668 ();
 sg13g2_fill_8 FILLER_0_71_676 ();
 sg13g2_fill_4 FILLER_0_71_684 ();
 sg13g2_fill_2 FILLER_0_71_688 ();
 sg13g2_fill_1 FILLER_0_71_690 ();
 sg13g2_fill_8 FILLER_0_71_696 ();
 sg13g2_fill_8 FILLER_0_71_704 ();
 sg13g2_fill_8 FILLER_0_71_712 ();
 sg13g2_fill_1 FILLER_0_71_720 ();
 sg13g2_fill_2 FILLER_0_71_731 ();
 sg13g2_fill_2 FILLER_0_71_739 ();
 sg13g2_fill_2 FILLER_0_71_751 ();
 sg13g2_fill_8 FILLER_0_71_779 ();
 sg13g2_fill_8 FILLER_0_71_787 ();
 sg13g2_fill_8 FILLER_0_71_795 ();
 sg13g2_fill_4 FILLER_0_71_803 ();
 sg13g2_fill_1 FILLER_0_71_807 ();
 sg13g2_fill_8 FILLER_0_71_813 ();
 sg13g2_fill_4 FILLER_0_71_826 ();
 sg13g2_fill_2 FILLER_0_71_830 ();
 sg13g2_fill_8 FILLER_0_71_837 ();
 sg13g2_fill_8 FILLER_0_71_845 ();
 sg13g2_fill_8 FILLER_0_71_853 ();
 sg13g2_fill_4 FILLER_0_71_861 ();
 sg13g2_fill_2 FILLER_0_71_865 ();
 sg13g2_fill_1 FILLER_0_71_867 ();
 sg13g2_fill_8 FILLER_0_71_873 ();
 sg13g2_fill_8 FILLER_0_71_881 ();
 sg13g2_fill_2 FILLER_0_71_889 ();
 sg13g2_fill_4 FILLER_0_71_896 ();
 sg13g2_fill_2 FILLER_0_71_900 ();
 sg13g2_fill_8 FILLER_0_71_912 ();
 sg13g2_fill_8 FILLER_0_71_926 ();
 sg13g2_fill_8 FILLER_0_71_934 ();
 sg13g2_fill_8 FILLER_0_71_946 ();
 sg13g2_fill_8 FILLER_0_71_954 ();
 sg13g2_fill_8 FILLER_0_71_962 ();
 sg13g2_fill_8 FILLER_0_71_975 ();
 sg13g2_fill_4 FILLER_0_71_983 ();
 sg13g2_fill_2 FILLER_0_71_987 ();
 sg13g2_fill_8 FILLER_0_71_994 ();
 sg13g2_fill_8 FILLER_0_71_1002 ();
 sg13g2_fill_4 FILLER_0_71_1010 ();
 sg13g2_fill_2 FILLER_0_71_1014 ();
 sg13g2_fill_8 FILLER_0_71_1020 ();
 sg13g2_fill_8 FILLER_0_71_1028 ();
 sg13g2_fill_2 FILLER_0_71_1036 ();
 sg13g2_fill_2 FILLER_0_71_1042 ();
 sg13g2_fill_1 FILLER_0_71_1044 ();
 sg13g2_fill_8 FILLER_0_71_1049 ();
 sg13g2_fill_8 FILLER_0_71_1063 ();
 sg13g2_fill_8 FILLER_0_71_1071 ();
 sg13g2_fill_4 FILLER_0_71_1079 ();
 sg13g2_fill_1 FILLER_0_71_1083 ();
 sg13g2_fill_8 FILLER_0_71_1088 ();
 sg13g2_fill_8 FILLER_0_71_1096 ();
 sg13g2_fill_2 FILLER_0_71_1104 ();
 sg13g2_fill_1 FILLER_0_71_1106 ();
 sg13g2_fill_2 FILLER_0_71_1111 ();
 sg13g2_fill_8 FILLER_0_71_1118 ();
 sg13g2_fill_8 FILLER_0_71_1126 ();
 sg13g2_fill_1 FILLER_0_71_1134 ();
 sg13g2_fill_4 FILLER_0_71_1139 ();
 sg13g2_fill_1 FILLER_0_71_1143 ();
 sg13g2_fill_2 FILLER_0_71_1148 ();
 sg13g2_fill_2 FILLER_0_71_1155 ();
 sg13g2_fill_4 FILLER_0_71_1161 ();
 sg13g2_fill_2 FILLER_0_71_1169 ();
 sg13g2_fill_1 FILLER_0_71_1171 ();
 sg13g2_fill_2 FILLER_0_71_1177 ();
 sg13g2_fill_4 FILLER_0_71_1184 ();
 sg13g2_fill_8 FILLER_0_71_1192 ();
 sg13g2_fill_8 FILLER_0_71_1200 ();
 sg13g2_fill_4 FILLER_0_71_1208 ();
 sg13g2_fill_2 FILLER_0_71_1212 ();
 sg13g2_fill_4 FILLER_0_71_1219 ();
 sg13g2_fill_2 FILLER_0_71_1231 ();
 sg13g2_fill_2 FILLER_0_71_1236 ();
 sg13g2_fill_2 FILLER_0_71_1242 ();
 sg13g2_fill_2 FILLER_0_71_1248 ();
 sg13g2_fill_1 FILLER_0_71_1250 ();
 sg13g2_fill_2 FILLER_0_71_1255 ();
 sg13g2_fill_1 FILLER_0_71_1257 ();
 sg13g2_fill_2 FILLER_0_71_1284 ();
 sg13g2_fill_4 FILLER_0_71_1290 ();
 sg13g2_fill_2 FILLER_0_71_1294 ();
 sg13g2_fill_1 FILLER_0_71_1296 ();
 sg13g2_fill_8 FILLER_0_72_0 ();
 sg13g2_fill_8 FILLER_0_72_8 ();
 sg13g2_fill_8 FILLER_0_72_16 ();
 sg13g2_fill_8 FILLER_0_72_24 ();
 sg13g2_fill_8 FILLER_0_72_32 ();
 sg13g2_fill_8 FILLER_0_72_40 ();
 sg13g2_fill_8 FILLER_0_72_48 ();
 sg13g2_fill_8 FILLER_0_72_56 ();
 sg13g2_fill_8 FILLER_0_72_64 ();
 sg13g2_fill_8 FILLER_0_72_72 ();
 sg13g2_fill_8 FILLER_0_72_80 ();
 sg13g2_fill_8 FILLER_0_72_88 ();
 sg13g2_fill_8 FILLER_0_72_96 ();
 sg13g2_fill_8 FILLER_0_72_104 ();
 sg13g2_fill_8 FILLER_0_72_112 ();
 sg13g2_fill_8 FILLER_0_72_120 ();
 sg13g2_fill_8 FILLER_0_72_128 ();
 sg13g2_fill_8 FILLER_0_72_136 ();
 sg13g2_fill_8 FILLER_0_72_144 ();
 sg13g2_fill_8 FILLER_0_72_152 ();
 sg13g2_fill_8 FILLER_0_72_160 ();
 sg13g2_fill_8 FILLER_0_72_168 ();
 sg13g2_fill_8 FILLER_0_72_176 ();
 sg13g2_fill_8 FILLER_0_72_184 ();
 sg13g2_fill_8 FILLER_0_72_192 ();
 sg13g2_fill_8 FILLER_0_72_200 ();
 sg13g2_fill_4 FILLER_0_72_208 ();
 sg13g2_fill_1 FILLER_0_72_212 ();
 sg13g2_fill_2 FILLER_0_72_218 ();
 sg13g2_fill_8 FILLER_0_72_246 ();
 sg13g2_fill_8 FILLER_0_72_260 ();
 sg13g2_fill_8 FILLER_0_72_268 ();
 sg13g2_fill_8 FILLER_0_72_276 ();
 sg13g2_fill_8 FILLER_0_72_284 ();
 sg13g2_fill_4 FILLER_0_72_292 ();
 sg13g2_fill_2 FILLER_0_72_296 ();
 sg13g2_fill_4 FILLER_0_72_302 ();
 sg13g2_fill_2 FILLER_0_72_311 ();
 sg13g2_fill_4 FILLER_0_72_318 ();
 sg13g2_fill_2 FILLER_0_72_322 ();
 sg13g2_fill_1 FILLER_0_72_324 ();
 sg13g2_fill_4 FILLER_0_72_329 ();
 sg13g2_fill_2 FILLER_0_72_338 ();
 sg13g2_fill_8 FILLER_0_72_348 ();
 sg13g2_fill_2 FILLER_0_72_356 ();
 sg13g2_fill_1 FILLER_0_72_358 ();
 sg13g2_fill_4 FILLER_0_72_363 ();
 sg13g2_fill_2 FILLER_0_72_367 ();
 sg13g2_fill_1 FILLER_0_72_369 ();
 sg13g2_fill_2 FILLER_0_72_375 ();
 sg13g2_fill_8 FILLER_0_72_383 ();
 sg13g2_fill_8 FILLER_0_72_391 ();
 sg13g2_fill_4 FILLER_0_72_399 ();
 sg13g2_fill_2 FILLER_0_72_408 ();
 sg13g2_fill_1 FILLER_0_72_410 ();
 sg13g2_fill_2 FILLER_0_72_415 ();
 sg13g2_fill_2 FILLER_0_72_420 ();
 sg13g2_fill_2 FILLER_0_72_427 ();
 sg13g2_fill_2 FILLER_0_72_433 ();
 sg13g2_fill_4 FILLER_0_72_441 ();
 sg13g2_fill_8 FILLER_0_72_466 ();
 sg13g2_fill_1 FILLER_0_72_474 ();
 sg13g2_fill_2 FILLER_0_72_481 ();
 sg13g2_fill_1 FILLER_0_72_483 ();
 sg13g2_fill_8 FILLER_0_72_488 ();
 sg13g2_fill_2 FILLER_0_72_496 ();
 sg13g2_fill_8 FILLER_0_72_503 ();
 sg13g2_fill_2 FILLER_0_72_511 ();
 sg13g2_fill_1 FILLER_0_72_513 ();
 sg13g2_fill_8 FILLER_0_72_519 ();
 sg13g2_fill_2 FILLER_0_72_527 ();
 sg13g2_fill_1 FILLER_0_72_529 ();
 sg13g2_fill_4 FILLER_0_72_534 ();
 sg13g2_fill_1 FILLER_0_72_538 ();
 sg13g2_fill_2 FILLER_0_72_565 ();
 sg13g2_fill_2 FILLER_0_72_572 ();
 sg13g2_fill_4 FILLER_0_72_578 ();
 sg13g2_fill_2 FILLER_0_72_582 ();
 sg13g2_fill_2 FILLER_0_72_589 ();
 sg13g2_fill_4 FILLER_0_72_596 ();
 sg13g2_fill_1 FILLER_0_72_600 ();
 sg13g2_fill_8 FILLER_0_72_605 ();
 sg13g2_fill_8 FILLER_0_72_613 ();
 sg13g2_fill_8 FILLER_0_72_621 ();
 sg13g2_fill_8 FILLER_0_72_629 ();
 sg13g2_fill_8 FILLER_0_72_637 ();
 sg13g2_fill_8 FILLER_0_72_645 ();
 sg13g2_fill_4 FILLER_0_72_653 ();
 sg13g2_fill_2 FILLER_0_72_667 ();
 sg13g2_fill_8 FILLER_0_72_674 ();
 sg13g2_fill_2 FILLER_0_72_682 ();
 sg13g2_fill_2 FILLER_0_72_694 ();
 sg13g2_fill_1 FILLER_0_72_696 ();
 sg13g2_fill_4 FILLER_0_72_723 ();
 sg13g2_fill_2 FILLER_0_72_732 ();
 sg13g2_fill_1 FILLER_0_72_734 ();
 sg13g2_fill_4 FILLER_0_72_741 ();
 sg13g2_fill_2 FILLER_0_72_771 ();
 sg13g2_fill_4 FILLER_0_72_783 ();
 sg13g2_fill_1 FILLER_0_72_787 ();
 sg13g2_fill_2 FILLER_0_72_793 ();
 sg13g2_fill_4 FILLER_0_72_821 ();
 sg13g2_fill_8 FILLER_0_72_851 ();
 sg13g2_fill_2 FILLER_0_72_859 ();
 sg13g2_fill_1 FILLER_0_72_861 ();
 sg13g2_fill_8 FILLER_0_72_866 ();
 sg13g2_fill_2 FILLER_0_72_874 ();
 sg13g2_fill_2 FILLER_0_72_880 ();
 sg13g2_fill_2 FILLER_0_72_887 ();
 sg13g2_fill_8 FILLER_0_72_892 ();
 sg13g2_fill_8 FILLER_0_72_900 ();
 sg13g2_fill_4 FILLER_0_72_908 ();
 sg13g2_fill_2 FILLER_0_72_912 ();
 sg13g2_fill_1 FILLER_0_72_914 ();
 sg13g2_fill_8 FILLER_0_72_920 ();
 sg13g2_fill_8 FILLER_0_72_928 ();
 sg13g2_fill_8 FILLER_0_72_936 ();
 sg13g2_fill_8 FILLER_0_72_944 ();
 sg13g2_fill_4 FILLER_0_72_952 ();
 sg13g2_fill_2 FILLER_0_72_956 ();
 sg13g2_fill_2 FILLER_0_72_963 ();
 sg13g2_fill_2 FILLER_0_72_969 ();
 sg13g2_fill_8 FILLER_0_72_978 ();
 sg13g2_fill_8 FILLER_0_72_986 ();
 sg13g2_fill_8 FILLER_0_72_994 ();
 sg13g2_fill_4 FILLER_0_72_1002 ();
 sg13g2_fill_2 FILLER_0_72_1010 ();
 sg13g2_fill_2 FILLER_0_72_1017 ();
 sg13g2_fill_1 FILLER_0_72_1019 ();
 sg13g2_fill_2 FILLER_0_72_1024 ();
 sg13g2_fill_4 FILLER_0_72_1033 ();
 sg13g2_fill_1 FILLER_0_72_1037 ();
 sg13g2_fill_8 FILLER_0_72_1043 ();
 sg13g2_fill_4 FILLER_0_72_1051 ();
 sg13g2_fill_2 FILLER_0_72_1055 ();
 sg13g2_fill_1 FILLER_0_72_1057 ();
 sg13g2_fill_8 FILLER_0_72_1063 ();
 sg13g2_fill_8 FILLER_0_72_1071 ();
 sg13g2_fill_4 FILLER_0_72_1079 ();
 sg13g2_fill_2 FILLER_0_72_1091 ();
 sg13g2_fill_2 FILLER_0_72_1097 ();
 sg13g2_fill_1 FILLER_0_72_1099 ();
 sg13g2_fill_2 FILLER_0_72_1108 ();
 sg13g2_fill_8 FILLER_0_72_1118 ();
 sg13g2_fill_2 FILLER_0_72_1134 ();
 sg13g2_fill_2 FILLER_0_72_1142 ();
 sg13g2_fill_8 FILLER_0_72_1149 ();
 sg13g2_fill_4 FILLER_0_72_1157 ();
 sg13g2_fill_1 FILLER_0_72_1161 ();
 sg13g2_fill_2 FILLER_0_72_1170 ();
 sg13g2_fill_8 FILLER_0_72_1177 ();
 sg13g2_fill_8 FILLER_0_72_1185 ();
 sg13g2_fill_8 FILLER_0_72_1193 ();
 sg13g2_fill_8 FILLER_0_72_1201 ();
 sg13g2_fill_8 FILLER_0_72_1209 ();
 sg13g2_fill_4 FILLER_0_72_1217 ();
 sg13g2_fill_2 FILLER_0_72_1221 ();
 sg13g2_fill_2 FILLER_0_72_1231 ();
 sg13g2_fill_1 FILLER_0_72_1233 ();
 sg13g2_fill_2 FILLER_0_72_1239 ();
 sg13g2_fill_2 FILLER_0_72_1249 ();
 sg13g2_fill_8 FILLER_0_72_1261 ();
 sg13g2_fill_4 FILLER_0_72_1269 ();
 sg13g2_fill_1 FILLER_0_72_1273 ();
 sg13g2_fill_2 FILLER_0_72_1282 ();
 sg13g2_fill_1 FILLER_0_72_1284 ();
 sg13g2_fill_8 FILLER_0_72_1289 ();
 sg13g2_fill_8 FILLER_0_73_0 ();
 sg13g2_fill_8 FILLER_0_73_8 ();
 sg13g2_fill_8 FILLER_0_73_16 ();
 sg13g2_fill_8 FILLER_0_73_24 ();
 sg13g2_fill_8 FILLER_0_73_32 ();
 sg13g2_fill_8 FILLER_0_73_40 ();
 sg13g2_fill_8 FILLER_0_73_48 ();
 sg13g2_fill_8 FILLER_0_73_56 ();
 sg13g2_fill_8 FILLER_0_73_64 ();
 sg13g2_fill_8 FILLER_0_73_72 ();
 sg13g2_fill_8 FILLER_0_73_80 ();
 sg13g2_fill_8 FILLER_0_73_88 ();
 sg13g2_fill_8 FILLER_0_73_96 ();
 sg13g2_fill_8 FILLER_0_73_104 ();
 sg13g2_fill_8 FILLER_0_73_112 ();
 sg13g2_fill_8 FILLER_0_73_120 ();
 sg13g2_fill_8 FILLER_0_73_128 ();
 sg13g2_fill_8 FILLER_0_73_136 ();
 sg13g2_fill_8 FILLER_0_73_144 ();
 sg13g2_fill_8 FILLER_0_73_152 ();
 sg13g2_fill_8 FILLER_0_73_160 ();
 sg13g2_fill_8 FILLER_0_73_168 ();
 sg13g2_fill_8 FILLER_0_73_176 ();
 sg13g2_fill_8 FILLER_0_73_184 ();
 sg13g2_fill_8 FILLER_0_73_192 ();
 sg13g2_fill_8 FILLER_0_73_200 ();
 sg13g2_fill_8 FILLER_0_73_208 ();
 sg13g2_fill_8 FILLER_0_73_216 ();
 sg13g2_fill_8 FILLER_0_73_224 ();
 sg13g2_fill_4 FILLER_0_73_232 ();
 sg13g2_fill_2 FILLER_0_73_236 ();
 sg13g2_fill_8 FILLER_0_73_264 ();
 sg13g2_fill_8 FILLER_0_73_272 ();
 sg13g2_fill_8 FILLER_0_73_280 ();
 sg13g2_fill_8 FILLER_0_73_288 ();
 sg13g2_fill_8 FILLER_0_73_296 ();
 sg13g2_fill_8 FILLER_0_73_304 ();
 sg13g2_fill_8 FILLER_0_73_312 ();
 sg13g2_fill_8 FILLER_0_73_320 ();
 sg13g2_fill_8 FILLER_0_73_328 ();
 sg13g2_fill_8 FILLER_0_73_336 ();
 sg13g2_fill_8 FILLER_0_73_344 ();
 sg13g2_fill_8 FILLER_0_73_352 ();
 sg13g2_fill_8 FILLER_0_73_360 ();
 sg13g2_fill_8 FILLER_0_73_368 ();
 sg13g2_fill_8 FILLER_0_73_376 ();
 sg13g2_fill_8 FILLER_0_73_384 ();
 sg13g2_fill_8 FILLER_0_73_392 ();
 sg13g2_fill_8 FILLER_0_73_400 ();
 sg13g2_fill_8 FILLER_0_73_408 ();
 sg13g2_fill_2 FILLER_0_73_416 ();
 sg13g2_fill_1 FILLER_0_73_418 ();
 sg13g2_fill_8 FILLER_0_73_425 ();
 sg13g2_fill_4 FILLER_0_73_433 ();
 sg13g2_fill_1 FILLER_0_73_437 ();
 sg13g2_fill_8 FILLER_0_73_443 ();
 sg13g2_fill_8 FILLER_0_73_451 ();
 sg13g2_fill_4 FILLER_0_73_459 ();
 sg13g2_fill_2 FILLER_0_73_467 ();
 sg13g2_fill_1 FILLER_0_73_469 ();
 sg13g2_fill_8 FILLER_0_73_476 ();
 sg13g2_fill_8 FILLER_0_73_484 ();
 sg13g2_fill_8 FILLER_0_73_492 ();
 sg13g2_fill_8 FILLER_0_73_500 ();
 sg13g2_fill_8 FILLER_0_73_508 ();
 sg13g2_fill_4 FILLER_0_73_516 ();
 sg13g2_fill_2 FILLER_0_73_520 ();
 sg13g2_fill_1 FILLER_0_73_522 ();
 sg13g2_fill_4 FILLER_0_73_528 ();
 sg13g2_fill_1 FILLER_0_73_532 ();
 sg13g2_fill_2 FILLER_0_73_537 ();
 sg13g2_fill_2 FILLER_0_73_565 ();
 sg13g2_fill_2 FILLER_0_73_572 ();
 sg13g2_fill_1 FILLER_0_73_574 ();
 sg13g2_fill_2 FILLER_0_73_579 ();
 sg13g2_fill_2 FILLER_0_73_607 ();
 sg13g2_fill_4 FILLER_0_73_630 ();
 sg13g2_fill_2 FILLER_0_73_634 ();
 sg13g2_fill_2 FILLER_0_73_662 ();
 sg13g2_fill_2 FILLER_0_73_669 ();
 sg13g2_fill_1 FILLER_0_73_671 ();
 sg13g2_fill_8 FILLER_0_73_682 ();
 sg13g2_fill_4 FILLER_0_73_690 ();
 sg13g2_fill_2 FILLER_0_73_694 ();
 sg13g2_fill_1 FILLER_0_73_696 ();
 sg13g2_fill_8 FILLER_0_73_723 ();
 sg13g2_fill_2 FILLER_0_73_731 ();
 sg13g2_fill_8 FILLER_0_73_738 ();
 sg13g2_fill_8 FILLER_0_73_746 ();
 sg13g2_fill_8 FILLER_0_73_754 ();
 sg13g2_fill_8 FILLER_0_73_762 ();
 sg13g2_fill_8 FILLER_0_73_770 ();
 sg13g2_fill_8 FILLER_0_73_778 ();
 sg13g2_fill_4 FILLER_0_73_786 ();
 sg13g2_fill_2 FILLER_0_73_790 ();
 sg13g2_fill_2 FILLER_0_73_797 ();
 sg13g2_fill_8 FILLER_0_73_809 ();
 sg13g2_fill_4 FILLER_0_73_817 ();
 sg13g2_fill_2 FILLER_0_73_826 ();
 sg13g2_fill_2 FILLER_0_73_833 ();
 sg13g2_fill_2 FILLER_0_73_845 ();
 sg13g2_fill_1 FILLER_0_73_847 ();
 sg13g2_fill_8 FILLER_0_73_853 ();
 sg13g2_fill_2 FILLER_0_73_861 ();
 sg13g2_fill_8 FILLER_0_73_867 ();
 sg13g2_fill_8 FILLER_0_73_875 ();
 sg13g2_fill_4 FILLER_0_73_883 ();
 sg13g2_fill_4 FILLER_0_73_892 ();
 sg13g2_fill_1 FILLER_0_73_896 ();
 sg13g2_fill_2 FILLER_0_73_902 ();
 sg13g2_fill_8 FILLER_0_73_925 ();
 sg13g2_fill_4 FILLER_0_73_933 ();
 sg13g2_fill_2 FILLER_0_73_937 ();
 sg13g2_fill_1 FILLER_0_73_939 ();
 sg13g2_fill_8 FILLER_0_73_945 ();
 sg13g2_fill_4 FILLER_0_73_953 ();
 sg13g2_fill_2 FILLER_0_73_957 ();
 sg13g2_fill_1 FILLER_0_73_959 ();
 sg13g2_fill_8 FILLER_0_73_965 ();
 sg13g2_fill_2 FILLER_0_73_977 ();
 sg13g2_fill_1 FILLER_0_73_979 ();
 sg13g2_fill_2 FILLER_0_73_985 ();
 sg13g2_fill_8 FILLER_0_73_993 ();
 sg13g2_fill_4 FILLER_0_73_1001 ();
 sg13g2_fill_1 FILLER_0_73_1005 ();
 sg13g2_fill_2 FILLER_0_73_1016 ();
 sg13g2_fill_2 FILLER_0_73_1023 ();
 sg13g2_fill_2 FILLER_0_73_1029 ();
 sg13g2_fill_8 FILLER_0_73_1036 ();
 sg13g2_fill_2 FILLER_0_73_1044 ();
 sg13g2_fill_8 FILLER_0_73_1051 ();
 sg13g2_fill_4 FILLER_0_73_1059 ();
 sg13g2_fill_1 FILLER_0_73_1063 ();
 sg13g2_fill_2 FILLER_0_73_1069 ();
 sg13g2_fill_8 FILLER_0_73_1077 ();
 sg13g2_fill_2 FILLER_0_73_1085 ();
 sg13g2_fill_1 FILLER_0_73_1087 ();
 sg13g2_fill_2 FILLER_0_73_1093 ();
 sg13g2_fill_2 FILLER_0_73_1100 ();
 sg13g2_fill_8 FILLER_0_73_1107 ();
 sg13g2_fill_4 FILLER_0_73_1115 ();
 sg13g2_fill_1 FILLER_0_73_1119 ();
 sg13g2_fill_4 FILLER_0_73_1124 ();
 sg13g2_fill_1 FILLER_0_73_1128 ();
 sg13g2_fill_2 FILLER_0_73_1134 ();
 sg13g2_fill_2 FILLER_0_73_1142 ();
 sg13g2_fill_8 FILLER_0_73_1149 ();
 sg13g2_fill_4 FILLER_0_73_1157 ();
 sg13g2_fill_1 FILLER_0_73_1161 ();
 sg13g2_fill_8 FILLER_0_73_1168 ();
 sg13g2_fill_4 FILLER_0_73_1176 ();
 sg13g2_fill_8 FILLER_0_73_1187 ();
 sg13g2_fill_8 FILLER_0_73_1195 ();
 sg13g2_fill_8 FILLER_0_73_1203 ();
 sg13g2_fill_4 FILLER_0_73_1211 ();
 sg13g2_fill_4 FILLER_0_73_1220 ();
 sg13g2_fill_1 FILLER_0_73_1224 ();
 sg13g2_fill_4 FILLER_0_73_1230 ();
 sg13g2_fill_2 FILLER_0_73_1234 ();
 sg13g2_fill_1 FILLER_0_73_1236 ();
 sg13g2_fill_8 FILLER_0_73_1242 ();
 sg13g2_fill_2 FILLER_0_73_1250 ();
 sg13g2_fill_1 FILLER_0_73_1252 ();
 sg13g2_fill_4 FILLER_0_73_1257 ();
 sg13g2_fill_2 FILLER_0_73_1261 ();
 sg13g2_fill_2 FILLER_0_73_1268 ();
 sg13g2_fill_8 FILLER_0_73_1274 ();
 sg13g2_fill_8 FILLER_0_73_1282 ();
 sg13g2_fill_4 FILLER_0_73_1290 ();
 sg13g2_fill_2 FILLER_0_73_1294 ();
 sg13g2_fill_1 FILLER_0_73_1296 ();
 sg13g2_fill_8 FILLER_0_74_0 ();
 sg13g2_fill_8 FILLER_0_74_8 ();
 sg13g2_fill_8 FILLER_0_74_16 ();
 sg13g2_fill_8 FILLER_0_74_24 ();
 sg13g2_fill_8 FILLER_0_74_32 ();
 sg13g2_fill_8 FILLER_0_74_40 ();
 sg13g2_fill_8 FILLER_0_74_48 ();
 sg13g2_fill_8 FILLER_0_74_56 ();
 sg13g2_fill_8 FILLER_0_74_64 ();
 sg13g2_fill_8 FILLER_0_74_72 ();
 sg13g2_fill_8 FILLER_0_74_80 ();
 sg13g2_fill_8 FILLER_0_74_88 ();
 sg13g2_fill_8 FILLER_0_74_96 ();
 sg13g2_fill_8 FILLER_0_74_104 ();
 sg13g2_fill_8 FILLER_0_74_112 ();
 sg13g2_fill_8 FILLER_0_74_120 ();
 sg13g2_fill_8 FILLER_0_74_128 ();
 sg13g2_fill_8 FILLER_0_74_136 ();
 sg13g2_fill_8 FILLER_0_74_144 ();
 sg13g2_fill_8 FILLER_0_74_152 ();
 sg13g2_fill_8 FILLER_0_74_160 ();
 sg13g2_fill_8 FILLER_0_74_168 ();
 sg13g2_fill_8 FILLER_0_74_176 ();
 sg13g2_fill_8 FILLER_0_74_184 ();
 sg13g2_fill_8 FILLER_0_74_192 ();
 sg13g2_fill_8 FILLER_0_74_200 ();
 sg13g2_fill_8 FILLER_0_74_208 ();
 sg13g2_fill_8 FILLER_0_74_216 ();
 sg13g2_fill_8 FILLER_0_74_224 ();
 sg13g2_fill_8 FILLER_0_74_232 ();
 sg13g2_fill_8 FILLER_0_74_240 ();
 sg13g2_fill_1 FILLER_0_74_248 ();
 sg13g2_fill_8 FILLER_0_74_254 ();
 sg13g2_fill_8 FILLER_0_74_262 ();
 sg13g2_fill_2 FILLER_0_74_270 ();
 sg13g2_fill_2 FILLER_0_74_277 ();
 sg13g2_fill_1 FILLER_0_74_279 ();
 sg13g2_fill_8 FILLER_0_74_284 ();
 sg13g2_fill_4 FILLER_0_74_292 ();
 sg13g2_fill_1 FILLER_0_74_296 ();
 sg13g2_fill_8 FILLER_0_74_318 ();
 sg13g2_fill_4 FILLER_0_74_326 ();
 sg13g2_fill_2 FILLER_0_74_330 ();
 sg13g2_fill_8 FILLER_0_74_336 ();
 sg13g2_fill_8 FILLER_0_74_344 ();
 sg13g2_fill_2 FILLER_0_74_356 ();
 sg13g2_fill_4 FILLER_0_74_362 ();
 sg13g2_fill_2 FILLER_0_74_366 ();
 sg13g2_fill_2 FILLER_0_74_389 ();
 sg13g2_fill_2 FILLER_0_74_396 ();
 sg13g2_fill_1 FILLER_0_74_398 ();
 sg13g2_fill_2 FILLER_0_74_403 ();
 sg13g2_fill_4 FILLER_0_74_410 ();
 sg13g2_fill_2 FILLER_0_74_414 ();
 sg13g2_fill_8 FILLER_0_74_421 ();
 sg13g2_fill_8 FILLER_0_74_429 ();
 sg13g2_fill_8 FILLER_0_74_437 ();
 sg13g2_fill_8 FILLER_0_74_445 ();
 sg13g2_fill_8 FILLER_0_74_453 ();
 sg13g2_fill_8 FILLER_0_74_461 ();
 sg13g2_fill_8 FILLER_0_74_469 ();
 sg13g2_fill_8 FILLER_0_74_477 ();
 sg13g2_fill_8 FILLER_0_74_485 ();
 sg13g2_fill_8 FILLER_0_74_493 ();
 sg13g2_fill_2 FILLER_0_74_501 ();
 sg13g2_fill_8 FILLER_0_74_515 ();
 sg13g2_fill_2 FILLER_0_74_530 ();
 sg13g2_fill_4 FILLER_0_74_537 ();
 sg13g2_fill_2 FILLER_0_74_546 ();
 sg13g2_fill_1 FILLER_0_74_548 ();
 sg13g2_fill_2 FILLER_0_74_554 ();
 sg13g2_fill_1 FILLER_0_74_556 ();
 sg13g2_fill_8 FILLER_0_74_567 ();
 sg13g2_fill_8 FILLER_0_74_575 ();
 sg13g2_fill_4 FILLER_0_74_588 ();
 sg13g2_fill_1 FILLER_0_74_592 ();
 sg13g2_fill_2 FILLER_0_74_619 ();
 sg13g2_fill_8 FILLER_0_74_625 ();
 sg13g2_fill_2 FILLER_0_74_633 ();
 sg13g2_fill_1 FILLER_0_74_635 ();
 sg13g2_fill_2 FILLER_0_74_662 ();
 sg13g2_fill_1 FILLER_0_74_664 ();
 sg13g2_fill_8 FILLER_0_74_691 ();
 sg13g2_fill_8 FILLER_0_74_699 ();
 sg13g2_fill_2 FILLER_0_74_712 ();
 sg13g2_fill_8 FILLER_0_74_719 ();
 sg13g2_fill_8 FILLER_0_74_727 ();
 sg13g2_fill_8 FILLER_0_74_735 ();
 sg13g2_fill_4 FILLER_0_74_743 ();
 sg13g2_fill_2 FILLER_0_74_747 ();
 sg13g2_fill_8 FILLER_0_74_759 ();
 sg13g2_fill_2 FILLER_0_74_767 ();
 sg13g2_fill_1 FILLER_0_74_769 ();
 sg13g2_fill_8 FILLER_0_74_791 ();
 sg13g2_fill_8 FILLER_0_74_799 ();
 sg13g2_fill_4 FILLER_0_74_807 ();
 sg13g2_fill_2 FILLER_0_74_811 ();
 sg13g2_fill_2 FILLER_0_74_817 ();
 sg13g2_fill_8 FILLER_0_74_823 ();
 sg13g2_fill_8 FILLER_0_74_831 ();
 sg13g2_fill_8 FILLER_0_74_839 ();
 sg13g2_fill_8 FILLER_0_74_847 ();
 sg13g2_fill_4 FILLER_0_74_855 ();
 sg13g2_fill_1 FILLER_0_74_859 ();
 sg13g2_fill_8 FILLER_0_74_864 ();
 sg13g2_fill_8 FILLER_0_74_872 ();
 sg13g2_fill_4 FILLER_0_74_885 ();
 sg13g2_fill_2 FILLER_0_74_889 ();
 sg13g2_fill_1 FILLER_0_74_891 ();
 sg13g2_fill_8 FILLER_0_74_902 ();
 sg13g2_fill_8 FILLER_0_74_910 ();
 sg13g2_fill_2 FILLER_0_74_918 ();
 sg13g2_fill_1 FILLER_0_74_920 ();
 sg13g2_fill_2 FILLER_0_74_925 ();
 sg13g2_fill_2 FILLER_0_74_933 ();
 sg13g2_fill_4 FILLER_0_74_939 ();
 sg13g2_fill_2 FILLER_0_74_943 ();
 sg13g2_fill_1 FILLER_0_74_945 ();
 sg13g2_fill_2 FILLER_0_74_953 ();
 sg13g2_fill_2 FILLER_0_74_960 ();
 sg13g2_fill_2 FILLER_0_74_966 ();
 sg13g2_fill_2 FILLER_0_74_978 ();
 sg13g2_fill_2 FILLER_0_74_988 ();
 sg13g2_fill_4 FILLER_0_74_994 ();
 sg13g2_fill_4 FILLER_0_74_1002 ();
 sg13g2_fill_8 FILLER_0_74_1016 ();
 sg13g2_fill_1 FILLER_0_74_1024 ();
 sg13g2_fill_2 FILLER_0_74_1029 ();
 sg13g2_fill_4 FILLER_0_74_1036 ();
 sg13g2_fill_2 FILLER_0_74_1040 ();
 sg13g2_fill_4 FILLER_0_74_1047 ();
 sg13g2_fill_4 FILLER_0_74_1056 ();
 sg13g2_fill_1 FILLER_0_74_1060 ();
 sg13g2_fill_4 FILLER_0_74_1066 ();
 sg13g2_fill_1 FILLER_0_74_1070 ();
 sg13g2_fill_4 FILLER_0_74_1078 ();
 sg13g2_fill_1 FILLER_0_74_1082 ();
 sg13g2_fill_4 FILLER_0_74_1088 ();
 sg13g2_fill_1 FILLER_0_74_1092 ();
 sg13g2_fill_2 FILLER_0_74_1098 ();
 sg13g2_fill_2 FILLER_0_74_1105 ();
 sg13g2_fill_2 FILLER_0_74_1112 ();
 sg13g2_fill_1 FILLER_0_74_1114 ();
 sg13g2_fill_8 FILLER_0_74_1120 ();
 sg13g2_fill_4 FILLER_0_74_1128 ();
 sg13g2_fill_2 FILLER_0_74_1132 ();
 sg13g2_fill_2 FILLER_0_74_1140 ();
 sg13g2_fill_2 FILLER_0_74_1147 ();
 sg13g2_fill_4 FILLER_0_74_1154 ();
 sg13g2_fill_2 FILLER_0_74_1164 ();
 sg13g2_fill_2 FILLER_0_74_1170 ();
 sg13g2_fill_2 FILLER_0_74_1177 ();
 sg13g2_fill_8 FILLER_0_74_1184 ();
 sg13g2_fill_8 FILLER_0_74_1192 ();
 sg13g2_fill_8 FILLER_0_74_1200 ();
 sg13g2_fill_1 FILLER_0_74_1208 ();
 sg13g2_fill_2 FILLER_0_74_1213 ();
 sg13g2_fill_2 FILLER_0_74_1220 ();
 sg13g2_fill_2 FILLER_0_74_1227 ();
 sg13g2_fill_8 FILLER_0_74_1234 ();
 sg13g2_fill_2 FILLER_0_74_1242 ();
 sg13g2_fill_1 FILLER_0_74_1244 ();
 sg13g2_fill_8 FILLER_0_74_1249 ();
 sg13g2_fill_8 FILLER_0_74_1262 ();
 sg13g2_fill_8 FILLER_0_74_1270 ();
 sg13g2_fill_2 FILLER_0_74_1278 ();
 sg13g2_fill_8 FILLER_0_74_1284 ();
 sg13g2_fill_4 FILLER_0_74_1292 ();
 sg13g2_fill_1 FILLER_0_74_1296 ();
 sg13g2_fill_8 FILLER_0_75_0 ();
 sg13g2_fill_8 FILLER_0_75_8 ();
 sg13g2_fill_8 FILLER_0_75_16 ();
 sg13g2_fill_8 FILLER_0_75_24 ();
 sg13g2_fill_8 FILLER_0_75_32 ();
 sg13g2_fill_8 FILLER_0_75_40 ();
 sg13g2_fill_8 FILLER_0_75_48 ();
 sg13g2_fill_8 FILLER_0_75_56 ();
 sg13g2_fill_8 FILLER_0_75_64 ();
 sg13g2_fill_8 FILLER_0_75_72 ();
 sg13g2_fill_8 FILLER_0_75_80 ();
 sg13g2_fill_8 FILLER_0_75_88 ();
 sg13g2_fill_8 FILLER_0_75_96 ();
 sg13g2_fill_8 FILLER_0_75_104 ();
 sg13g2_fill_8 FILLER_0_75_112 ();
 sg13g2_fill_8 FILLER_0_75_120 ();
 sg13g2_fill_8 FILLER_0_75_128 ();
 sg13g2_fill_8 FILLER_0_75_136 ();
 sg13g2_fill_8 FILLER_0_75_144 ();
 sg13g2_fill_8 FILLER_0_75_152 ();
 sg13g2_fill_8 FILLER_0_75_160 ();
 sg13g2_fill_8 FILLER_0_75_168 ();
 sg13g2_fill_8 FILLER_0_75_176 ();
 sg13g2_fill_8 FILLER_0_75_184 ();
 sg13g2_fill_8 FILLER_0_75_192 ();
 sg13g2_fill_8 FILLER_0_75_200 ();
 sg13g2_fill_8 FILLER_0_75_208 ();
 sg13g2_fill_8 FILLER_0_75_216 ();
 sg13g2_fill_8 FILLER_0_75_224 ();
 sg13g2_fill_8 FILLER_0_75_232 ();
 sg13g2_fill_8 FILLER_0_75_240 ();
 sg13g2_fill_8 FILLER_0_75_248 ();
 sg13g2_fill_8 FILLER_0_75_256 ();
 sg13g2_fill_4 FILLER_0_75_264 ();
 sg13g2_fill_1 FILLER_0_75_268 ();
 sg13g2_fill_2 FILLER_0_75_295 ();
 sg13g2_fill_2 FILLER_0_75_301 ();
 sg13g2_fill_1 FILLER_0_75_303 ();
 sg13g2_fill_2 FILLER_0_75_330 ();
 sg13g2_fill_8 FILLER_0_75_337 ();
 sg13g2_fill_2 FILLER_0_75_371 ();
 sg13g2_fill_2 FILLER_0_75_378 ();
 sg13g2_fill_8 FILLER_0_75_385 ();
 sg13g2_fill_8 FILLER_0_75_393 ();
 sg13g2_fill_1 FILLER_0_75_401 ();
 sg13g2_fill_8 FILLER_0_75_407 ();
 sg13g2_fill_2 FILLER_0_75_415 ();
 sg13g2_fill_2 FILLER_0_75_443 ();
 sg13g2_fill_1 FILLER_0_75_445 ();
 sg13g2_fill_2 FILLER_0_75_452 ();
 sg13g2_fill_2 FILLER_0_75_460 ();
 sg13g2_fill_2 FILLER_0_75_467 ();
 sg13g2_fill_2 FILLER_0_75_473 ();
 sg13g2_fill_2 FILLER_0_75_479 ();
 sg13g2_fill_8 FILLER_0_75_507 ();
 sg13g2_fill_8 FILLER_0_75_515 ();
 sg13g2_fill_2 FILLER_0_75_530 ();
 sg13g2_fill_8 FILLER_0_75_537 ();
 sg13g2_fill_8 FILLER_0_75_545 ();
 sg13g2_fill_1 FILLER_0_75_553 ();
 sg13g2_fill_8 FILLER_0_75_559 ();
 sg13g2_fill_8 FILLER_0_75_567 ();
 sg13g2_fill_8 FILLER_0_75_575 ();
 sg13g2_fill_8 FILLER_0_75_583 ();
 sg13g2_fill_1 FILLER_0_75_591 ();
 sg13g2_fill_2 FILLER_0_75_597 ();
 sg13g2_fill_8 FILLER_0_75_609 ();
 sg13g2_fill_8 FILLER_0_75_617 ();
 sg13g2_fill_8 FILLER_0_75_625 ();
 sg13g2_fill_4 FILLER_0_75_633 ();
 sg13g2_fill_2 FILLER_0_75_637 ();
 sg13g2_fill_2 FILLER_0_75_649 ();
 sg13g2_fill_1 FILLER_0_75_651 ();
 sg13g2_fill_2 FILLER_0_75_673 ();
 sg13g2_fill_1 FILLER_0_75_675 ();
 sg13g2_fill_8 FILLER_0_75_686 ();
 sg13g2_fill_4 FILLER_0_75_694 ();
 sg13g2_fill_1 FILLER_0_75_698 ();
 sg13g2_fill_8 FILLER_0_75_704 ();
 sg13g2_fill_1 FILLER_0_75_712 ();
 sg13g2_fill_4 FILLER_0_75_717 ();
 sg13g2_fill_1 FILLER_0_75_721 ();
 sg13g2_fill_8 FILLER_0_75_726 ();
 sg13g2_fill_8 FILLER_0_75_734 ();
 sg13g2_fill_8 FILLER_0_75_742 ();
 sg13g2_fill_4 FILLER_0_75_750 ();
 sg13g2_fill_2 FILLER_0_75_754 ();
 sg13g2_fill_1 FILLER_0_75_756 ();
 sg13g2_fill_8 FILLER_0_75_783 ();
 sg13g2_fill_8 FILLER_0_75_791 ();
 sg13g2_fill_4 FILLER_0_75_799 ();
 sg13g2_fill_8 FILLER_0_75_807 ();
 sg13g2_fill_8 FILLER_0_75_815 ();
 sg13g2_fill_8 FILLER_0_75_823 ();
 sg13g2_fill_8 FILLER_0_75_831 ();
 sg13g2_fill_8 FILLER_0_75_839 ();
 sg13g2_fill_8 FILLER_0_75_847 ();
 sg13g2_fill_8 FILLER_0_75_855 ();
 sg13g2_fill_8 FILLER_0_75_863 ();
 sg13g2_fill_8 FILLER_0_75_871 ();
 sg13g2_fill_8 FILLER_0_75_879 ();
 sg13g2_fill_2 FILLER_0_75_887 ();
 sg13g2_fill_2 FILLER_0_75_893 ();
 sg13g2_fill_1 FILLER_0_75_895 ();
 sg13g2_fill_8 FILLER_0_75_906 ();
 sg13g2_fill_2 FILLER_0_75_914 ();
 sg13g2_fill_4 FILLER_0_75_920 ();
 sg13g2_fill_4 FILLER_0_75_929 ();
 sg13g2_fill_8 FILLER_0_75_939 ();
 sg13g2_fill_8 FILLER_0_75_947 ();
 sg13g2_fill_4 FILLER_0_75_955 ();
 sg13g2_fill_2 FILLER_0_75_965 ();
 sg13g2_fill_2 FILLER_0_75_972 ();
 sg13g2_fill_4 FILLER_0_75_978 ();
 sg13g2_fill_2 FILLER_0_75_982 ();
 sg13g2_fill_1 FILLER_0_75_984 ();
 sg13g2_fill_8 FILLER_0_75_990 ();
 sg13g2_fill_8 FILLER_0_75_998 ();
 sg13g2_fill_8 FILLER_0_75_1006 ();
 sg13g2_fill_8 FILLER_0_75_1014 ();
 sg13g2_fill_4 FILLER_0_75_1022 ();
 sg13g2_fill_8 FILLER_0_75_1031 ();
 sg13g2_fill_2 FILLER_0_75_1039 ();
 sg13g2_fill_8 FILLER_0_75_1045 ();
 sg13g2_fill_8 FILLER_0_75_1053 ();
 sg13g2_fill_8 FILLER_0_75_1061 ();
 sg13g2_fill_8 FILLER_0_75_1069 ();
 sg13g2_fill_4 FILLER_0_75_1077 ();
 sg13g2_fill_8 FILLER_0_75_1086 ();
 sg13g2_fill_2 FILLER_0_75_1094 ();
 sg13g2_fill_8 FILLER_0_75_1101 ();
 sg13g2_fill_4 FILLER_0_75_1109 ();
 sg13g2_fill_8 FILLER_0_75_1122 ();
 sg13g2_fill_4 FILLER_0_75_1130 ();
 sg13g2_fill_4 FILLER_0_75_1140 ();
 sg13g2_fill_2 FILLER_0_75_1150 ();
 sg13g2_fill_1 FILLER_0_75_1152 ();
 sg13g2_fill_4 FILLER_0_75_1158 ();
 sg13g2_fill_1 FILLER_0_75_1162 ();
 sg13g2_fill_2 FILLER_0_75_1167 ();
 sg13g2_fill_2 FILLER_0_75_1174 ();
 sg13g2_fill_2 FILLER_0_75_1184 ();
 sg13g2_fill_4 FILLER_0_75_1194 ();
 sg13g2_fill_1 FILLER_0_75_1198 ();
 sg13g2_fill_8 FILLER_0_75_1204 ();
 sg13g2_fill_1 FILLER_0_75_1212 ();
 sg13g2_fill_2 FILLER_0_75_1219 ();
 sg13g2_fill_8 FILLER_0_75_1226 ();
 sg13g2_fill_8 FILLER_0_75_1239 ();
 sg13g2_fill_4 FILLER_0_75_1247 ();
 sg13g2_fill_1 FILLER_0_75_1251 ();
 sg13g2_fill_2 FILLER_0_75_1256 ();
 sg13g2_fill_2 FILLER_0_75_1284 ();
 sg13g2_fill_2 FILLER_0_75_1290 ();
 sg13g2_fill_1 FILLER_0_75_1296 ();
 sg13g2_fill_8 FILLER_0_76_0 ();
 sg13g2_fill_8 FILLER_0_76_8 ();
 sg13g2_fill_8 FILLER_0_76_16 ();
 sg13g2_fill_8 FILLER_0_76_24 ();
 sg13g2_fill_8 FILLER_0_76_32 ();
 sg13g2_fill_8 FILLER_0_76_40 ();
 sg13g2_fill_8 FILLER_0_76_48 ();
 sg13g2_fill_8 FILLER_0_76_56 ();
 sg13g2_fill_8 FILLER_0_76_64 ();
 sg13g2_fill_8 FILLER_0_76_72 ();
 sg13g2_fill_8 FILLER_0_76_80 ();
 sg13g2_fill_8 FILLER_0_76_88 ();
 sg13g2_fill_8 FILLER_0_76_96 ();
 sg13g2_fill_8 FILLER_0_76_104 ();
 sg13g2_fill_8 FILLER_0_76_112 ();
 sg13g2_fill_8 FILLER_0_76_120 ();
 sg13g2_fill_8 FILLER_0_76_128 ();
 sg13g2_fill_8 FILLER_0_76_136 ();
 sg13g2_fill_8 FILLER_0_76_144 ();
 sg13g2_fill_8 FILLER_0_76_152 ();
 sg13g2_fill_8 FILLER_0_76_160 ();
 sg13g2_fill_8 FILLER_0_76_168 ();
 sg13g2_fill_8 FILLER_0_76_176 ();
 sg13g2_fill_8 FILLER_0_76_184 ();
 sg13g2_fill_8 FILLER_0_76_192 ();
 sg13g2_fill_8 FILLER_0_76_200 ();
 sg13g2_fill_8 FILLER_0_76_208 ();
 sg13g2_fill_4 FILLER_0_76_216 ();
 sg13g2_fill_2 FILLER_0_76_220 ();
 sg13g2_fill_1 FILLER_0_76_222 ();
 sg13g2_fill_8 FILLER_0_76_249 ();
 sg13g2_fill_8 FILLER_0_76_257 ();
 sg13g2_fill_4 FILLER_0_76_265 ();
 sg13g2_fill_1 FILLER_0_76_269 ();
 sg13g2_fill_4 FILLER_0_76_296 ();
 sg13g2_fill_1 FILLER_0_76_300 ();
 sg13g2_fill_8 FILLER_0_76_322 ();
 sg13g2_fill_8 FILLER_0_76_330 ();
 sg13g2_fill_4 FILLER_0_76_338 ();
 sg13g2_fill_2 FILLER_0_76_342 ();
 sg13g2_fill_1 FILLER_0_76_344 ();
 sg13g2_fill_2 FILLER_0_76_371 ();
 sg13g2_fill_1 FILLER_0_76_373 ();
 sg13g2_fill_4 FILLER_0_76_379 ();
 sg13g2_fill_2 FILLER_0_76_383 ();
 sg13g2_fill_2 FILLER_0_76_390 ();
 sg13g2_fill_2 FILLER_0_76_397 ();
 sg13g2_fill_4 FILLER_0_76_404 ();
 sg13g2_fill_2 FILLER_0_76_408 ();
 sg13g2_fill_1 FILLER_0_76_410 ();
 sg13g2_fill_4 FILLER_0_76_416 ();
 sg13g2_fill_2 FILLER_0_76_420 ();
 sg13g2_fill_1 FILLER_0_76_422 ();
 sg13g2_fill_2 FILLER_0_76_428 ();
 sg13g2_fill_8 FILLER_0_76_434 ();
 sg13g2_fill_8 FILLER_0_76_448 ();
 sg13g2_fill_2 FILLER_0_76_466 ();
 sg13g2_fill_2 FILLER_0_76_473 ();
 sg13g2_fill_2 FILLER_0_76_480 ();
 sg13g2_fill_2 FILLER_0_76_508 ();
 sg13g2_fill_8 FILLER_0_76_520 ();
 sg13g2_fill_2 FILLER_0_76_528 ();
 sg13g2_fill_1 FILLER_0_76_530 ();
 sg13g2_fill_2 FILLER_0_76_537 ();
 sg13g2_fill_1 FILLER_0_76_539 ();
 sg13g2_fill_4 FILLER_0_76_545 ();
 sg13g2_fill_1 FILLER_0_76_549 ();
 sg13g2_fill_2 FILLER_0_76_556 ();
 sg13g2_fill_8 FILLER_0_76_563 ();
 sg13g2_fill_8 FILLER_0_76_571 ();
 sg13g2_fill_1 FILLER_0_76_579 ();
 sg13g2_fill_8 FILLER_0_76_588 ();
 sg13g2_fill_8 FILLER_0_76_596 ();
 sg13g2_fill_8 FILLER_0_76_604 ();
 sg13g2_fill_8 FILLER_0_76_612 ();
 sg13g2_fill_8 FILLER_0_76_620 ();
 sg13g2_fill_8 FILLER_0_76_628 ();
 sg13g2_fill_8 FILLER_0_76_636 ();
 sg13g2_fill_8 FILLER_0_76_644 ();
 sg13g2_fill_4 FILLER_0_76_652 ();
 sg13g2_fill_2 FILLER_0_76_656 ();
 sg13g2_fill_4 FILLER_0_76_668 ();
 sg13g2_fill_2 FILLER_0_76_672 ();
 sg13g2_fill_8 FILLER_0_76_678 ();
 sg13g2_fill_2 FILLER_0_76_691 ();
 sg13g2_fill_4 FILLER_0_76_701 ();
 sg13g2_fill_2 FILLER_0_76_705 ();
 sg13g2_fill_2 FILLER_0_76_711 ();
 sg13g2_fill_4 FILLER_0_76_734 ();
 sg13g2_fill_2 FILLER_0_76_738 ();
 sg13g2_fill_1 FILLER_0_76_740 ();
 sg13g2_fill_2 FILLER_0_76_751 ();
 sg13g2_fill_4 FILLER_0_76_779 ();
 sg13g2_fill_4 FILLER_0_76_791 ();
 sg13g2_fill_8 FILLER_0_76_821 ();
 sg13g2_fill_8 FILLER_0_76_855 ();
 sg13g2_fill_8 FILLER_0_76_863 ();
 sg13g2_fill_8 FILLER_0_76_871 ();
 sg13g2_fill_2 FILLER_0_76_879 ();
 sg13g2_fill_1 FILLER_0_76_881 ();
 sg13g2_fill_2 FILLER_0_76_886 ();
 sg13g2_fill_8 FILLER_0_76_893 ();
 sg13g2_fill_4 FILLER_0_76_901 ();
 sg13g2_fill_8 FILLER_0_76_926 ();
 sg13g2_fill_8 FILLER_0_76_934 ();
 sg13g2_fill_8 FILLER_0_76_942 ();
 sg13g2_fill_8 FILLER_0_76_950 ();
 sg13g2_fill_4 FILLER_0_76_958 ();
 sg13g2_fill_2 FILLER_0_76_962 ();
 sg13g2_fill_8 FILLER_0_76_969 ();
 sg13g2_fill_8 FILLER_0_76_982 ();
 sg13g2_fill_8 FILLER_0_76_990 ();
 sg13g2_fill_8 FILLER_0_76_998 ();
 sg13g2_fill_8 FILLER_0_76_1006 ();
 sg13g2_fill_4 FILLER_0_76_1014 ();
 sg13g2_fill_8 FILLER_0_76_1023 ();
 sg13g2_fill_1 FILLER_0_76_1031 ();
 sg13g2_fill_8 FILLER_0_76_1038 ();
 sg13g2_fill_1 FILLER_0_76_1046 ();
 sg13g2_fill_8 FILLER_0_76_1052 ();
 sg13g2_fill_8 FILLER_0_76_1060 ();
 sg13g2_fill_8 FILLER_0_76_1068 ();
 sg13g2_fill_8 FILLER_0_76_1076 ();
 sg13g2_fill_8 FILLER_0_76_1084 ();
 sg13g2_fill_8 FILLER_0_76_1092 ();
 sg13g2_fill_8 FILLER_0_76_1100 ();
 sg13g2_fill_8 FILLER_0_76_1108 ();
 sg13g2_fill_2 FILLER_0_76_1120 ();
 sg13g2_fill_8 FILLER_0_76_1127 ();
 sg13g2_fill_4 FILLER_0_76_1140 ();
 sg13g2_fill_4 FILLER_0_76_1147 ();
 sg13g2_fill_2 FILLER_0_76_1151 ();
 sg13g2_fill_8 FILLER_0_76_1159 ();
 sg13g2_fill_2 FILLER_0_76_1167 ();
 sg13g2_fill_8 FILLER_0_76_1179 ();
 sg13g2_fill_8 FILLER_0_76_1187 ();
 sg13g2_fill_8 FILLER_0_76_1195 ();
 sg13g2_fill_8 FILLER_0_76_1203 ();
 sg13g2_fill_8 FILLER_0_76_1211 ();
 sg13g2_fill_1 FILLER_0_76_1219 ();
 sg13g2_fill_2 FILLER_0_76_1224 ();
 sg13g2_fill_2 FILLER_0_76_1230 ();
 sg13g2_fill_8 FILLER_0_76_1240 ();
 sg13g2_fill_1 FILLER_0_76_1248 ();
 sg13g2_fill_8 FILLER_0_76_1259 ();
 sg13g2_fill_8 FILLER_0_76_1267 ();
 sg13g2_fill_8 FILLER_0_76_1275 ();
 sg13g2_fill_8 FILLER_0_76_1283 ();
 sg13g2_fill_1 FILLER_0_76_1291 ();
 sg13g2_fill_1 FILLER_0_76_1296 ();
 sg13g2_fill_8 FILLER_0_77_0 ();
 sg13g2_fill_8 FILLER_0_77_8 ();
 sg13g2_fill_8 FILLER_0_77_16 ();
 sg13g2_fill_8 FILLER_0_77_24 ();
 sg13g2_fill_8 FILLER_0_77_32 ();
 sg13g2_fill_8 FILLER_0_77_40 ();
 sg13g2_fill_8 FILLER_0_77_48 ();
 sg13g2_fill_8 FILLER_0_77_56 ();
 sg13g2_fill_8 FILLER_0_77_64 ();
 sg13g2_fill_8 FILLER_0_77_72 ();
 sg13g2_fill_8 FILLER_0_77_80 ();
 sg13g2_fill_8 FILLER_0_77_88 ();
 sg13g2_fill_8 FILLER_0_77_96 ();
 sg13g2_fill_8 FILLER_0_77_104 ();
 sg13g2_fill_8 FILLER_0_77_112 ();
 sg13g2_fill_8 FILLER_0_77_120 ();
 sg13g2_fill_8 FILLER_0_77_128 ();
 sg13g2_fill_8 FILLER_0_77_136 ();
 sg13g2_fill_8 FILLER_0_77_144 ();
 sg13g2_fill_8 FILLER_0_77_152 ();
 sg13g2_fill_8 FILLER_0_77_160 ();
 sg13g2_fill_8 FILLER_0_77_168 ();
 sg13g2_fill_8 FILLER_0_77_176 ();
 sg13g2_fill_8 FILLER_0_77_184 ();
 sg13g2_fill_8 FILLER_0_77_192 ();
 sg13g2_fill_8 FILLER_0_77_200 ();
 sg13g2_fill_8 FILLER_0_77_208 ();
 sg13g2_fill_8 FILLER_0_77_216 ();
 sg13g2_fill_4 FILLER_0_77_224 ();
 sg13g2_fill_2 FILLER_0_77_228 ();
 sg13g2_fill_8 FILLER_0_77_235 ();
 sg13g2_fill_1 FILLER_0_77_243 ();
 sg13g2_fill_8 FILLER_0_77_248 ();
 sg13g2_fill_2 FILLER_0_77_256 ();
 sg13g2_fill_2 FILLER_0_77_263 ();
 sg13g2_fill_2 FILLER_0_77_270 ();
 sg13g2_fill_2 FILLER_0_77_277 ();
 sg13g2_fill_8 FILLER_0_77_305 ();
 sg13g2_fill_8 FILLER_0_77_313 ();
 sg13g2_fill_8 FILLER_0_77_321 ();
 sg13g2_fill_8 FILLER_0_77_329 ();
 sg13g2_fill_2 FILLER_0_77_337 ();
 sg13g2_fill_1 FILLER_0_77_339 ();
 sg13g2_fill_4 FILLER_0_77_345 ();
 sg13g2_fill_1 FILLER_0_77_349 ();
 sg13g2_fill_2 FILLER_0_77_355 ();
 sg13g2_fill_4 FILLER_0_77_361 ();
 sg13g2_fill_2 FILLER_0_77_365 ();
 sg13g2_fill_4 FILLER_0_77_372 ();
 sg13g2_fill_2 FILLER_0_77_376 ();
 sg13g2_fill_1 FILLER_0_77_378 ();
 sg13g2_fill_2 FILLER_0_77_383 ();
 sg13g2_fill_4 FILLER_0_77_391 ();
 sg13g2_fill_8 FILLER_0_77_421 ();
 sg13g2_fill_1 FILLER_0_77_429 ();
 sg13g2_fill_8 FILLER_0_77_435 ();
 sg13g2_fill_4 FILLER_0_77_443 ();
 sg13g2_fill_1 FILLER_0_77_447 ();
 sg13g2_fill_8 FILLER_0_77_453 ();
 sg13g2_fill_8 FILLER_0_77_461 ();
 sg13g2_fill_8 FILLER_0_77_469 ();
 sg13g2_fill_4 FILLER_0_77_477 ();
 sg13g2_fill_1 FILLER_0_77_481 ();
 sg13g2_fill_8 FILLER_0_77_486 ();
 sg13g2_fill_4 FILLER_0_77_494 ();
 sg13g2_fill_8 FILLER_0_77_503 ();
 sg13g2_fill_8 FILLER_0_77_511 ();
 sg13g2_fill_4 FILLER_0_77_519 ();
 sg13g2_fill_1 FILLER_0_77_523 ();
 sg13g2_fill_8 FILLER_0_77_529 ();
 sg13g2_fill_2 FILLER_0_77_537 ();
 sg13g2_fill_8 FILLER_0_77_565 ();
 sg13g2_fill_8 FILLER_0_77_573 ();
 sg13g2_fill_4 FILLER_0_77_581 ();
 sg13g2_fill_8 FILLER_0_77_589 ();
 sg13g2_fill_1 FILLER_0_77_597 ();
 sg13g2_fill_2 FILLER_0_77_603 ();
 sg13g2_fill_8 FILLER_0_77_610 ();
 sg13g2_fill_8 FILLER_0_77_618 ();
 sg13g2_fill_8 FILLER_0_77_626 ();
 sg13g2_fill_8 FILLER_0_77_634 ();
 sg13g2_fill_2 FILLER_0_77_642 ();
 sg13g2_fill_1 FILLER_0_77_644 ();
 sg13g2_fill_8 FILLER_0_77_671 ();
 sg13g2_fill_2 FILLER_0_77_684 ();
 sg13g2_fill_8 FILLER_0_77_692 ();
 sg13g2_fill_4 FILLER_0_77_700 ();
 sg13g2_fill_1 FILLER_0_77_704 ();
 sg13g2_fill_2 FILLER_0_77_731 ();
 sg13g2_fill_4 FILLER_0_77_737 ();
 sg13g2_fill_4 FILLER_0_77_762 ();
 sg13g2_fill_1 FILLER_0_77_766 ();
 sg13g2_fill_2 FILLER_0_77_779 ();
 sg13g2_fill_1 FILLER_0_77_781 ();
 sg13g2_fill_2 FILLER_0_77_787 ();
 sg13g2_fill_1 FILLER_0_77_789 ();
 sg13g2_fill_4 FILLER_0_77_800 ();
 sg13g2_fill_2 FILLER_0_77_830 ();
 sg13g2_fill_8 FILLER_0_77_842 ();
 sg13g2_fill_2 FILLER_0_77_850 ();
 sg13g2_fill_1 FILLER_0_77_852 ();
 sg13g2_fill_8 FILLER_0_77_858 ();
 sg13g2_fill_8 FILLER_0_77_866 ();
 sg13g2_fill_8 FILLER_0_77_874 ();
 sg13g2_fill_4 FILLER_0_77_882 ();
 sg13g2_fill_2 FILLER_0_77_891 ();
 sg13g2_fill_8 FILLER_0_77_903 ();
 sg13g2_fill_8 FILLER_0_77_911 ();
 sg13g2_fill_4 FILLER_0_77_919 ();
 sg13g2_fill_1 FILLER_0_77_923 ();
 sg13g2_fill_2 FILLER_0_77_929 ();
 sg13g2_fill_4 FILLER_0_77_941 ();
 sg13g2_fill_2 FILLER_0_77_945 ();
 sg13g2_fill_8 FILLER_0_77_951 ();
 sg13g2_fill_1 FILLER_0_77_959 ();
 sg13g2_fill_2 FILLER_0_77_964 ();
 sg13g2_fill_8 FILLER_0_77_971 ();
 sg13g2_fill_2 FILLER_0_77_984 ();
 sg13g2_fill_8 FILLER_0_77_991 ();
 sg13g2_fill_4 FILLER_0_77_999 ();
 sg13g2_fill_2 FILLER_0_77_1003 ();
 sg13g2_fill_4 FILLER_0_77_1011 ();
 sg13g2_fill_2 FILLER_0_77_1023 ();
 sg13g2_fill_1 FILLER_0_77_1025 ();
 sg13g2_fill_2 FILLER_0_77_1032 ();
 sg13g2_fill_2 FILLER_0_77_1038 ();
 sg13g2_fill_4 FILLER_0_77_1044 ();
 sg13g2_fill_2 FILLER_0_77_1053 ();
 sg13g2_fill_8 FILLER_0_77_1062 ();
 sg13g2_fill_8 FILLER_0_77_1070 ();
 sg13g2_fill_8 FILLER_0_77_1078 ();
 sg13g2_fill_8 FILLER_0_77_1086 ();
 sg13g2_fill_8 FILLER_0_77_1094 ();
 sg13g2_fill_8 FILLER_0_77_1102 ();
 sg13g2_fill_4 FILLER_0_77_1110 ();
 sg13g2_fill_2 FILLER_0_77_1114 ();
 sg13g2_fill_1 FILLER_0_77_1116 ();
 sg13g2_fill_8 FILLER_0_77_1122 ();
 sg13g2_fill_2 FILLER_0_77_1134 ();
 sg13g2_fill_8 FILLER_0_77_1139 ();
 sg13g2_fill_8 FILLER_0_77_1147 ();
 sg13g2_fill_8 FILLER_0_77_1155 ();
 sg13g2_fill_8 FILLER_0_77_1163 ();
 sg13g2_fill_4 FILLER_0_77_1171 ();
 sg13g2_fill_2 FILLER_0_77_1175 ();
 sg13g2_fill_8 FILLER_0_77_1182 ();
 sg13g2_fill_8 FILLER_0_77_1190 ();
 sg13g2_fill_8 FILLER_0_77_1198 ();
 sg13g2_fill_8 FILLER_0_77_1206 ();
 sg13g2_fill_8 FILLER_0_77_1214 ();
 sg13g2_fill_8 FILLER_0_77_1222 ();
 sg13g2_fill_8 FILLER_0_77_1230 ();
 sg13g2_fill_4 FILLER_0_77_1238 ();
 sg13g2_fill_2 FILLER_0_77_1242 ();
 sg13g2_fill_2 FILLER_0_77_1254 ();
 sg13g2_fill_8 FILLER_0_77_1261 ();
 sg13g2_fill_8 FILLER_0_77_1269 ();
 sg13g2_fill_2 FILLER_0_77_1277 ();
 sg13g2_fill_8 FILLER_0_77_1287 ();
 sg13g2_fill_2 FILLER_0_77_1295 ();
 sg13g2_fill_8 FILLER_0_78_0 ();
 sg13g2_fill_8 FILLER_0_78_8 ();
 sg13g2_fill_8 FILLER_0_78_16 ();
 sg13g2_fill_8 FILLER_0_78_24 ();
 sg13g2_fill_8 FILLER_0_78_32 ();
 sg13g2_fill_8 FILLER_0_78_40 ();
 sg13g2_fill_8 FILLER_0_78_48 ();
 sg13g2_fill_8 FILLER_0_78_56 ();
 sg13g2_fill_8 FILLER_0_78_64 ();
 sg13g2_fill_8 FILLER_0_78_72 ();
 sg13g2_fill_8 FILLER_0_78_80 ();
 sg13g2_fill_8 FILLER_0_78_88 ();
 sg13g2_fill_8 FILLER_0_78_96 ();
 sg13g2_fill_8 FILLER_0_78_104 ();
 sg13g2_fill_8 FILLER_0_78_112 ();
 sg13g2_fill_8 FILLER_0_78_120 ();
 sg13g2_fill_8 FILLER_0_78_128 ();
 sg13g2_fill_8 FILLER_0_78_136 ();
 sg13g2_fill_8 FILLER_0_78_144 ();
 sg13g2_fill_8 FILLER_0_78_152 ();
 sg13g2_fill_8 FILLER_0_78_160 ();
 sg13g2_fill_8 FILLER_0_78_168 ();
 sg13g2_fill_8 FILLER_0_78_176 ();
 sg13g2_fill_8 FILLER_0_78_184 ();
 sg13g2_fill_8 FILLER_0_78_192 ();
 sg13g2_fill_8 FILLER_0_78_200 ();
 sg13g2_fill_8 FILLER_0_78_213 ();
 sg13g2_fill_4 FILLER_0_78_225 ();
 sg13g2_fill_2 FILLER_0_78_229 ();
 sg13g2_fill_1 FILLER_0_78_231 ();
 sg13g2_fill_2 FILLER_0_78_258 ();
 sg13g2_fill_8 FILLER_0_78_264 ();
 sg13g2_fill_8 FILLER_0_78_272 ();
 sg13g2_fill_2 FILLER_0_78_280 ();
 sg13g2_fill_2 FILLER_0_78_287 ();
 sg13g2_fill_1 FILLER_0_78_289 ();
 sg13g2_fill_8 FILLER_0_78_294 ();
 sg13g2_fill_8 FILLER_0_78_302 ();
 sg13g2_fill_8 FILLER_0_78_310 ();
 sg13g2_fill_8 FILLER_0_78_318 ();
 sg13g2_fill_8 FILLER_0_78_326 ();
 sg13g2_fill_8 FILLER_0_78_334 ();
 sg13g2_fill_8 FILLER_0_78_342 ();
 sg13g2_fill_8 FILLER_0_78_350 ();
 sg13g2_fill_8 FILLER_0_78_358 ();
 sg13g2_fill_8 FILLER_0_78_366 ();
 sg13g2_fill_8 FILLER_0_78_374 ();
 sg13g2_fill_8 FILLER_0_78_382 ();
 sg13g2_fill_8 FILLER_0_78_390 ();
 sg13g2_fill_8 FILLER_0_78_398 ();
 sg13g2_fill_2 FILLER_0_78_410 ();
 sg13g2_fill_1 FILLER_0_78_412 ();
 sg13g2_fill_8 FILLER_0_78_418 ();
 sg13g2_fill_8 FILLER_0_78_426 ();
 sg13g2_fill_4 FILLER_0_78_434 ();
 sg13g2_fill_1 FILLER_0_78_438 ();
 sg13g2_fill_4 FILLER_0_78_444 ();
 sg13g2_fill_2 FILLER_0_78_448 ();
 sg13g2_fill_1 FILLER_0_78_450 ();
 sg13g2_fill_2 FILLER_0_78_455 ();
 sg13g2_fill_1 FILLER_0_78_457 ();
 sg13g2_fill_8 FILLER_0_78_462 ();
 sg13g2_fill_1 FILLER_0_78_470 ();
 sg13g2_fill_8 FILLER_0_78_475 ();
 sg13g2_fill_8 FILLER_0_78_483 ();
 sg13g2_fill_8 FILLER_0_78_491 ();
 sg13g2_fill_8 FILLER_0_78_499 ();
 sg13g2_fill_8 FILLER_0_78_507 ();
 sg13g2_fill_2 FILLER_0_78_515 ();
 sg13g2_fill_1 FILLER_0_78_517 ();
 sg13g2_fill_8 FILLER_0_78_523 ();
 sg13g2_fill_8 FILLER_0_78_531 ();
 sg13g2_fill_4 FILLER_0_78_544 ();
 sg13g2_fill_2 FILLER_0_78_548 ();
 sg13g2_fill_8 FILLER_0_78_554 ();
 sg13g2_fill_8 FILLER_0_78_562 ();
 sg13g2_fill_8 FILLER_0_78_570 ();
 sg13g2_fill_2 FILLER_0_78_604 ();
 sg13g2_fill_8 FILLER_0_78_611 ();
 sg13g2_fill_8 FILLER_0_78_619 ();
 sg13g2_fill_8 FILLER_0_78_627 ();
 sg13g2_fill_2 FILLER_0_78_635 ();
 sg13g2_fill_1 FILLER_0_78_637 ();
 sg13g2_fill_8 FILLER_0_78_648 ();
 sg13g2_fill_8 FILLER_0_78_656 ();
 sg13g2_fill_8 FILLER_0_78_664 ();
 sg13g2_fill_8 FILLER_0_78_672 ();
 sg13g2_fill_2 FILLER_0_78_685 ();
 sg13g2_fill_8 FILLER_0_78_692 ();
 sg13g2_fill_8 FILLER_0_78_700 ();
 sg13g2_fill_4 FILLER_0_78_708 ();
 sg13g2_fill_1 FILLER_0_78_712 ();
 sg13g2_fill_2 FILLER_0_78_719 ();
 sg13g2_fill_2 FILLER_0_78_731 ();
 sg13g2_fill_8 FILLER_0_78_738 ();
 sg13g2_fill_8 FILLER_0_78_746 ();
 sg13g2_fill_8 FILLER_0_78_754 ();
 sg13g2_fill_2 FILLER_0_78_762 ();
 sg13g2_fill_8 FILLER_0_78_769 ();
 sg13g2_fill_8 FILLER_0_78_777 ();
 sg13g2_fill_8 FILLER_0_78_785 ();
 sg13g2_fill_8 FILLER_0_78_793 ();
 sg13g2_fill_2 FILLER_0_78_801 ();
 sg13g2_fill_1 FILLER_0_78_803 ();
 sg13g2_fill_2 FILLER_0_78_814 ();
 sg13g2_fill_2 FILLER_0_78_837 ();
 sg13g2_fill_2 FILLER_0_78_865 ();
 sg13g2_fill_4 FILLER_0_78_872 ();
 sg13g2_fill_2 FILLER_0_78_876 ();
 sg13g2_fill_2 FILLER_0_78_883 ();
 sg13g2_fill_2 FILLER_0_78_895 ();
 sg13g2_fill_1 FILLER_0_78_897 ();
 sg13g2_fill_4 FILLER_0_78_902 ();
 sg13g2_fill_2 FILLER_0_78_906 ();
 sg13g2_fill_2 FILLER_0_78_913 ();
 sg13g2_fill_2 FILLER_0_78_920 ();
 sg13g2_fill_4 FILLER_0_78_926 ();
 sg13g2_fill_2 FILLER_0_78_930 ();
 sg13g2_fill_1 FILLER_0_78_932 ();
 sg13g2_fill_2 FILLER_0_78_943 ();
 sg13g2_fill_1 FILLER_0_78_945 ();
 sg13g2_fill_2 FILLER_0_78_951 ();
 sg13g2_fill_8 FILLER_0_78_958 ();
 sg13g2_fill_8 FILLER_0_78_966 ();
 sg13g2_fill_4 FILLER_0_78_974 ();
 sg13g2_fill_2 FILLER_0_78_985 ();
 sg13g2_fill_8 FILLER_0_78_995 ();
 sg13g2_fill_4 FILLER_0_78_1003 ();
 sg13g2_fill_4 FILLER_0_78_1013 ();
 sg13g2_fill_2 FILLER_0_78_1023 ();
 sg13g2_fill_2 FILLER_0_78_1030 ();
 sg13g2_fill_1 FILLER_0_78_1032 ();
 sg13g2_fill_2 FILLER_0_78_1038 ();
 sg13g2_fill_2 FILLER_0_78_1045 ();
 sg13g2_fill_1 FILLER_0_78_1047 ();
 sg13g2_fill_4 FILLER_0_78_1053 ();
 sg13g2_fill_2 FILLER_0_78_1063 ();
 sg13g2_fill_8 FILLER_0_78_1070 ();
 sg13g2_fill_8 FILLER_0_78_1078 ();
 sg13g2_fill_8 FILLER_0_78_1086 ();
 sg13g2_fill_4 FILLER_0_78_1094 ();
 sg13g2_fill_2 FILLER_0_78_1108 ();
 sg13g2_fill_2 FILLER_0_78_1118 ();
 sg13g2_fill_1 FILLER_0_78_1120 ();
 sg13g2_fill_2 FILLER_0_78_1128 ();
 sg13g2_fill_2 FILLER_0_78_1134 ();
 sg13g2_fill_8 FILLER_0_78_1144 ();
 sg13g2_fill_2 FILLER_0_78_1156 ();
 sg13g2_fill_2 FILLER_0_78_1164 ();
 sg13g2_fill_8 FILLER_0_78_1171 ();
 sg13g2_fill_2 FILLER_0_78_1179 ();
 sg13g2_fill_1 FILLER_0_78_1181 ();
 sg13g2_fill_2 FILLER_0_78_1186 ();
 sg13g2_fill_8 FILLER_0_78_1196 ();
 sg13g2_fill_4 FILLER_0_78_1209 ();
 sg13g2_fill_2 FILLER_0_78_1221 ();
 sg13g2_fill_8 FILLER_0_78_1228 ();
 sg13g2_fill_2 FILLER_0_78_1241 ();
 sg13g2_fill_8 FILLER_0_78_1248 ();
 sg13g2_fill_4 FILLER_0_78_1256 ();
 sg13g2_fill_1 FILLER_0_78_1260 ();
 sg13g2_fill_8 FILLER_0_78_1267 ();
 sg13g2_fill_1 FILLER_0_78_1275 ();
 sg13g2_fill_2 FILLER_0_78_1280 ();
 sg13g2_fill_4 FILLER_0_78_1286 ();
 sg13g2_fill_2 FILLER_0_78_1290 ();
 sg13g2_fill_1 FILLER_0_78_1296 ();
 sg13g2_fill_8 FILLER_0_79_0 ();
 sg13g2_fill_8 FILLER_0_79_8 ();
 sg13g2_fill_8 FILLER_0_79_16 ();
 sg13g2_fill_8 FILLER_0_79_24 ();
 sg13g2_fill_8 FILLER_0_79_32 ();
 sg13g2_fill_8 FILLER_0_79_40 ();
 sg13g2_fill_8 FILLER_0_79_48 ();
 sg13g2_fill_8 FILLER_0_79_56 ();
 sg13g2_fill_8 FILLER_0_79_64 ();
 sg13g2_fill_8 FILLER_0_79_72 ();
 sg13g2_fill_8 FILLER_0_79_80 ();
 sg13g2_fill_8 FILLER_0_79_88 ();
 sg13g2_fill_8 FILLER_0_79_96 ();
 sg13g2_fill_8 FILLER_0_79_104 ();
 sg13g2_fill_8 FILLER_0_79_112 ();
 sg13g2_fill_8 FILLER_0_79_120 ();
 sg13g2_fill_8 FILLER_0_79_128 ();
 sg13g2_fill_8 FILLER_0_79_136 ();
 sg13g2_fill_8 FILLER_0_79_144 ();
 sg13g2_fill_8 FILLER_0_79_152 ();
 sg13g2_fill_8 FILLER_0_79_160 ();
 sg13g2_fill_8 FILLER_0_79_168 ();
 sg13g2_fill_8 FILLER_0_79_176 ();
 sg13g2_fill_8 FILLER_0_79_184 ();
 sg13g2_fill_8 FILLER_0_79_192 ();
 sg13g2_fill_2 FILLER_0_79_200 ();
 sg13g2_fill_1 FILLER_0_79_202 ();
 sg13g2_fill_8 FILLER_0_79_229 ();
 sg13g2_fill_8 FILLER_0_79_237 ();
 sg13g2_fill_8 FILLER_0_79_245 ();
 sg13g2_fill_1 FILLER_0_79_253 ();
 sg13g2_fill_8 FILLER_0_79_275 ();
 sg13g2_fill_8 FILLER_0_79_283 ();
 sg13g2_fill_8 FILLER_0_79_291 ();
 sg13g2_fill_8 FILLER_0_79_299 ();
 sg13g2_fill_8 FILLER_0_79_307 ();
 sg13g2_fill_8 FILLER_0_79_315 ();
 sg13g2_fill_4 FILLER_0_79_323 ();
 sg13g2_fill_1 FILLER_0_79_327 ();
 sg13g2_fill_2 FILLER_0_79_333 ();
 sg13g2_fill_8 FILLER_0_79_339 ();
 sg13g2_fill_8 FILLER_0_79_347 ();
 sg13g2_fill_8 FILLER_0_79_355 ();
 sg13g2_fill_4 FILLER_0_79_363 ();
 sg13g2_fill_2 FILLER_0_79_367 ();
 sg13g2_fill_8 FILLER_0_79_373 ();
 sg13g2_fill_4 FILLER_0_79_381 ();
 sg13g2_fill_1 FILLER_0_79_385 ();
 sg13g2_fill_2 FILLER_0_79_391 ();
 sg13g2_fill_8 FILLER_0_79_397 ();
 sg13g2_fill_8 FILLER_0_79_405 ();
 sg13g2_fill_8 FILLER_0_79_413 ();
 sg13g2_fill_8 FILLER_0_79_421 ();
 sg13g2_fill_4 FILLER_0_79_429 ();
 sg13g2_fill_2 FILLER_0_79_433 ();
 sg13g2_fill_1 FILLER_0_79_435 ();
 sg13g2_fill_8 FILLER_0_79_462 ();
 sg13g2_fill_8 FILLER_0_79_470 ();
 sg13g2_fill_4 FILLER_0_79_483 ();
 sg13g2_fill_1 FILLER_0_79_487 ();
 sg13g2_fill_8 FILLER_0_79_493 ();
 sg13g2_fill_8 FILLER_0_79_501 ();
 sg13g2_fill_8 FILLER_0_79_509 ();
 sg13g2_fill_8 FILLER_0_79_517 ();
 sg13g2_fill_4 FILLER_0_79_525 ();
 sg13g2_fill_8 FILLER_0_79_534 ();
 sg13g2_fill_4 FILLER_0_79_542 ();
 sg13g2_fill_2 FILLER_0_79_546 ();
 sg13g2_fill_2 FILLER_0_79_553 ();
 sg13g2_fill_8 FILLER_0_79_581 ();
 sg13g2_fill_8 FILLER_0_79_589 ();
 sg13g2_fill_4 FILLER_0_79_597 ();
 sg13g2_fill_2 FILLER_0_79_601 ();
 sg13g2_fill_8 FILLER_0_79_607 ();
 sg13g2_fill_8 FILLER_0_79_615 ();
 sg13g2_fill_8 FILLER_0_79_623 ();
 sg13g2_fill_8 FILLER_0_79_631 ();
 sg13g2_fill_8 FILLER_0_79_639 ();
 sg13g2_fill_8 FILLER_0_79_647 ();
 sg13g2_fill_1 FILLER_0_79_655 ();
 sg13g2_fill_2 FILLER_0_79_666 ();
 sg13g2_fill_2 FILLER_0_79_678 ();
 sg13g2_fill_2 FILLER_0_79_706 ();
 sg13g2_fill_2 FILLER_0_79_734 ();
 sg13g2_fill_2 FILLER_0_79_746 ();
 sg13g2_fill_1 FILLER_0_79_748 ();
 sg13g2_fill_8 FILLER_0_79_754 ();
 sg13g2_fill_8 FILLER_0_79_762 ();
 sg13g2_fill_8 FILLER_0_79_770 ();
 sg13g2_fill_8 FILLER_0_79_778 ();
 sg13g2_fill_8 FILLER_0_79_786 ();
 sg13g2_fill_4 FILLER_0_79_794 ();
 sg13g2_fill_2 FILLER_0_79_798 ();
 sg13g2_fill_1 FILLER_0_79_800 ();
 sg13g2_fill_2 FILLER_0_79_811 ();
 sg13g2_fill_2 FILLER_0_79_818 ();
 sg13g2_fill_4 FILLER_0_79_825 ();
 sg13g2_fill_1 FILLER_0_79_829 ();
 sg13g2_fill_8 FILLER_0_79_840 ();
 sg13g2_fill_8 FILLER_0_79_853 ();
 sg13g2_fill_4 FILLER_0_79_861 ();
 sg13g2_fill_2 FILLER_0_79_865 ();
 sg13g2_fill_1 FILLER_0_79_867 ();
 sg13g2_fill_8 FILLER_0_79_872 ();
 sg13g2_fill_8 FILLER_0_79_880 ();
 sg13g2_fill_8 FILLER_0_79_888 ();
 sg13g2_fill_8 FILLER_0_79_896 ();
 sg13g2_fill_8 FILLER_0_79_904 ();
 sg13g2_fill_4 FILLER_0_79_912 ();
 sg13g2_fill_1 FILLER_0_79_916 ();
 sg13g2_fill_4 FILLER_0_79_921 ();
 sg13g2_fill_4 FILLER_0_79_930 ();
 sg13g2_fill_2 FILLER_0_79_939 ();
 sg13g2_fill_2 FILLER_0_79_948 ();
 sg13g2_fill_8 FILLER_0_79_954 ();
 sg13g2_fill_2 FILLER_0_79_966 ();
 sg13g2_fill_2 FILLER_0_79_974 ();
 sg13g2_fill_4 FILLER_0_79_982 ();
 sg13g2_fill_1 FILLER_0_79_986 ();
 sg13g2_fill_8 FILLER_0_79_992 ();
 sg13g2_fill_8 FILLER_0_79_1000 ();
 sg13g2_fill_4 FILLER_0_79_1012 ();
 sg13g2_fill_2 FILLER_0_79_1022 ();
 sg13g2_fill_4 FILLER_0_79_1028 ();
 sg13g2_fill_1 FILLER_0_79_1032 ();
 sg13g2_fill_2 FILLER_0_79_1041 ();
 sg13g2_fill_4 FILLER_0_79_1048 ();
 sg13g2_fill_2 FILLER_0_79_1052 ();
 sg13g2_fill_2 FILLER_0_79_1059 ();
 sg13g2_fill_2 FILLER_0_79_1071 ();
 sg13g2_fill_2 FILLER_0_79_1078 ();
 sg13g2_fill_2 FILLER_0_79_1086 ();
 sg13g2_fill_8 FILLER_0_79_1093 ();
 sg13g2_fill_4 FILLER_0_79_1101 ();
 sg13g2_fill_2 FILLER_0_79_1105 ();
 sg13g2_fill_1 FILLER_0_79_1107 ();
 sg13g2_fill_4 FILLER_0_79_1112 ();
 sg13g2_fill_1 FILLER_0_79_1116 ();
 sg13g2_fill_2 FILLER_0_79_1122 ();
 sg13g2_fill_2 FILLER_0_79_1129 ();
 sg13g2_fill_2 FILLER_0_79_1139 ();
 sg13g2_fill_2 FILLER_0_79_1146 ();
 sg13g2_fill_1 FILLER_0_79_1148 ();
 sg13g2_fill_2 FILLER_0_79_1154 ();
 sg13g2_fill_2 FILLER_0_79_1163 ();
 sg13g2_fill_8 FILLER_0_79_1169 ();
 sg13g2_fill_8 FILLER_0_79_1177 ();
 sg13g2_fill_2 FILLER_0_79_1185 ();
 sg13g2_fill_2 FILLER_0_79_1192 ();
 sg13g2_fill_8 FILLER_0_79_1198 ();
 sg13g2_fill_4 FILLER_0_79_1206 ();
 sg13g2_fill_2 FILLER_0_79_1216 ();
 sg13g2_fill_1 FILLER_0_79_1218 ();
 sg13g2_fill_8 FILLER_0_79_1224 ();
 sg13g2_fill_2 FILLER_0_79_1236 ();
 sg13g2_fill_8 FILLER_0_79_1242 ();
 sg13g2_fill_4 FILLER_0_79_1250 ();
 sg13g2_fill_2 FILLER_0_79_1254 ();
 sg13g2_fill_2 FILLER_0_79_1260 ();
 sg13g2_fill_2 FILLER_0_79_1267 ();
 sg13g2_fill_8 FILLER_0_79_1274 ();
 sg13g2_fill_4 FILLER_0_79_1287 ();
 sg13g2_fill_1 FILLER_0_79_1291 ();
 sg13g2_fill_1 FILLER_0_79_1296 ();
 sg13g2_fill_8 FILLER_0_80_0 ();
 sg13g2_fill_8 FILLER_0_80_8 ();
 sg13g2_fill_8 FILLER_0_80_16 ();
 sg13g2_fill_8 FILLER_0_80_24 ();
 sg13g2_fill_8 FILLER_0_80_32 ();
 sg13g2_fill_8 FILLER_0_80_40 ();
 sg13g2_fill_8 FILLER_0_80_48 ();
 sg13g2_fill_8 FILLER_0_80_56 ();
 sg13g2_fill_8 FILLER_0_80_64 ();
 sg13g2_fill_8 FILLER_0_80_72 ();
 sg13g2_fill_8 FILLER_0_80_80 ();
 sg13g2_fill_8 FILLER_0_80_88 ();
 sg13g2_fill_8 FILLER_0_80_96 ();
 sg13g2_fill_8 FILLER_0_80_104 ();
 sg13g2_fill_8 FILLER_0_80_112 ();
 sg13g2_fill_8 FILLER_0_80_120 ();
 sg13g2_fill_8 FILLER_0_80_128 ();
 sg13g2_fill_8 FILLER_0_80_136 ();
 sg13g2_fill_8 FILLER_0_80_144 ();
 sg13g2_fill_8 FILLER_0_80_152 ();
 sg13g2_fill_8 FILLER_0_80_160 ();
 sg13g2_fill_8 FILLER_0_80_168 ();
 sg13g2_fill_8 FILLER_0_80_176 ();
 sg13g2_fill_8 FILLER_0_80_184 ();
 sg13g2_fill_8 FILLER_0_80_192 ();
 sg13g2_fill_4 FILLER_0_80_200 ();
 sg13g2_fill_2 FILLER_0_80_204 ();
 sg13g2_fill_8 FILLER_0_80_232 ();
 sg13g2_fill_4 FILLER_0_80_261 ();
 sg13g2_fill_2 FILLER_0_80_265 ();
 sg13g2_fill_2 FILLER_0_80_272 ();
 sg13g2_fill_2 FILLER_0_80_279 ();
 sg13g2_fill_2 FILLER_0_80_285 ();
 sg13g2_fill_2 FILLER_0_80_292 ();
 sg13g2_fill_8 FILLER_0_80_299 ();
 sg13g2_fill_8 FILLER_0_80_307 ();
 sg13g2_fill_4 FILLER_0_80_315 ();
 sg13g2_fill_2 FILLER_0_80_345 ();
 sg13g2_fill_2 FILLER_0_80_368 ();
 sg13g2_fill_4 FILLER_0_80_375 ();
 sg13g2_fill_2 FILLER_0_80_379 ();
 sg13g2_fill_1 FILLER_0_80_381 ();
 sg13g2_fill_8 FILLER_0_80_408 ();
 sg13g2_fill_8 FILLER_0_80_424 ();
 sg13g2_fill_2 FILLER_0_80_436 ();
 sg13g2_fill_4 FILLER_0_80_443 ();
 sg13g2_fill_2 FILLER_0_80_447 ();
 sg13g2_fill_1 FILLER_0_80_449 ();
 sg13g2_fill_8 FILLER_0_80_460 ();
 sg13g2_fill_8 FILLER_0_80_468 ();
 sg13g2_fill_4 FILLER_0_80_476 ();
 sg13g2_fill_8 FILLER_0_80_485 ();
 sg13g2_fill_4 FILLER_0_80_498 ();
 sg13g2_fill_2 FILLER_0_80_502 ();
 sg13g2_fill_4 FILLER_0_80_509 ();
 sg13g2_fill_2 FILLER_0_80_513 ();
 sg13g2_fill_1 FILLER_0_80_515 ();
 sg13g2_fill_2 FILLER_0_80_521 ();
 sg13g2_fill_1 FILLER_0_80_523 ();
 sg13g2_fill_8 FILLER_0_80_550 ();
 sg13g2_fill_2 FILLER_0_80_558 ();
 sg13g2_fill_4 FILLER_0_80_565 ();
 sg13g2_fill_8 FILLER_0_80_573 ();
 sg13g2_fill_1 FILLER_0_80_581 ();
 sg13g2_fill_2 FILLER_0_80_592 ();
 sg13g2_fill_2 FILLER_0_80_599 ();
 sg13g2_fill_2 FILLER_0_80_606 ();
 sg13g2_fill_4 FILLER_0_80_612 ();
 sg13g2_fill_2 FILLER_0_80_616 ();
 sg13g2_fill_2 FILLER_0_80_622 ();
 sg13g2_fill_8 FILLER_0_80_630 ();
 sg13g2_fill_8 FILLER_0_80_638 ();
 sg13g2_fill_8 FILLER_0_80_646 ();
 sg13g2_fill_4 FILLER_0_80_654 ();
 sg13g2_fill_2 FILLER_0_80_668 ();
 sg13g2_fill_4 FILLER_0_80_675 ();
 sg13g2_fill_4 FILLER_0_80_683 ();
 sg13g2_fill_1 FILLER_0_80_687 ();
 sg13g2_fill_4 FILLER_0_80_692 ();
 sg13g2_fill_2 FILLER_0_80_696 ();
 sg13g2_fill_4 FILLER_0_80_702 ();
 sg13g2_fill_2 FILLER_0_80_706 ();
 sg13g2_fill_8 FILLER_0_80_713 ();
 sg13g2_fill_8 FILLER_0_80_721 ();
 sg13g2_fill_8 FILLER_0_80_729 ();
 sg13g2_fill_8 FILLER_0_80_737 ();
 sg13g2_fill_8 FILLER_0_80_745 ();
 sg13g2_fill_2 FILLER_0_80_753 ();
 sg13g2_fill_2 FILLER_0_80_765 ();
 sg13g2_fill_1 FILLER_0_80_767 ();
 sg13g2_fill_2 FILLER_0_80_772 ();
 sg13g2_fill_8 FILLER_0_80_778 ();
 sg13g2_fill_8 FILLER_0_80_786 ();
 sg13g2_fill_8 FILLER_0_80_794 ();
 sg13g2_fill_4 FILLER_0_80_802 ();
 sg13g2_fill_2 FILLER_0_80_811 ();
 sg13g2_fill_2 FILLER_0_80_818 ();
 sg13g2_fill_2 FILLER_0_80_825 ();
 sg13g2_fill_2 FILLER_0_80_831 ();
 sg13g2_fill_8 FILLER_0_80_836 ();
 sg13g2_fill_8 FILLER_0_80_848 ();
 sg13g2_fill_8 FILLER_0_80_856 ();
 sg13g2_fill_8 FILLER_0_80_864 ();
 sg13g2_fill_8 FILLER_0_80_872 ();
 sg13g2_fill_8 FILLER_0_80_880 ();
 sg13g2_fill_4 FILLER_0_80_888 ();
 sg13g2_fill_2 FILLER_0_80_892 ();
 sg13g2_fill_8 FILLER_0_80_899 ();
 sg13g2_fill_8 FILLER_0_80_907 ();
 sg13g2_fill_4 FILLER_0_80_915 ();
 sg13g2_fill_2 FILLER_0_80_919 ();
 sg13g2_fill_2 FILLER_0_80_931 ();
 sg13g2_fill_4 FILLER_0_80_937 ();
 sg13g2_fill_1 FILLER_0_80_941 ();
 sg13g2_fill_4 FILLER_0_80_947 ();
 sg13g2_fill_1 FILLER_0_80_951 ();
 sg13g2_fill_4 FILLER_0_80_956 ();
 sg13g2_fill_1 FILLER_0_80_960 ();
 sg13g2_fill_4 FILLER_0_80_966 ();
 sg13g2_fill_1 FILLER_0_80_970 ();
 sg13g2_fill_2 FILLER_0_80_975 ();
 sg13g2_fill_8 FILLER_0_80_983 ();
 sg13g2_fill_8 FILLER_0_80_996 ();
 sg13g2_fill_4 FILLER_0_80_1004 ();
 sg13g2_fill_1 FILLER_0_80_1008 ();
 sg13g2_fill_2 FILLER_0_80_1015 ();
 sg13g2_fill_8 FILLER_0_80_1021 ();
 sg13g2_fill_8 FILLER_0_80_1029 ();
 sg13g2_fill_2 FILLER_0_80_1037 ();
 sg13g2_fill_1 FILLER_0_80_1039 ();
 sg13g2_fill_2 FILLER_0_80_1045 ();
 sg13g2_fill_8 FILLER_0_80_1053 ();
 sg13g2_fill_8 FILLER_0_80_1061 ();
 sg13g2_fill_8 FILLER_0_80_1069 ();
 sg13g2_fill_4 FILLER_0_80_1077 ();
 sg13g2_fill_8 FILLER_0_80_1086 ();
 sg13g2_fill_8 FILLER_0_80_1094 ();
 sg13g2_fill_8 FILLER_0_80_1102 ();
 sg13g2_fill_2 FILLER_0_80_1110 ();
 sg13g2_fill_1 FILLER_0_80_1112 ();
 sg13g2_fill_8 FILLER_0_80_1118 ();
 sg13g2_fill_8 FILLER_0_80_1126 ();
 sg13g2_fill_8 FILLER_0_80_1134 ();
 sg13g2_fill_2 FILLER_0_80_1142 ();
 sg13g2_fill_4 FILLER_0_80_1149 ();
 sg13g2_fill_2 FILLER_0_80_1153 ();
 sg13g2_fill_8 FILLER_0_80_1159 ();
 sg13g2_fill_2 FILLER_0_80_1167 ();
 sg13g2_fill_1 FILLER_0_80_1169 ();
 sg13g2_fill_8 FILLER_0_80_1174 ();
 sg13g2_fill_2 FILLER_0_80_1182 ();
 sg13g2_fill_1 FILLER_0_80_1184 ();
 sg13g2_fill_2 FILLER_0_80_1189 ();
 sg13g2_fill_2 FILLER_0_80_1195 ();
 sg13g2_fill_4 FILLER_0_80_1202 ();
 sg13g2_fill_1 FILLER_0_80_1206 ();
 sg13g2_fill_4 FILLER_0_80_1211 ();
 sg13g2_fill_1 FILLER_0_80_1215 ();
 sg13g2_fill_2 FILLER_0_80_1221 ();
 sg13g2_fill_2 FILLER_0_80_1227 ();
 sg13g2_fill_1 FILLER_0_80_1229 ();
 sg13g2_fill_8 FILLER_0_80_1238 ();
 sg13g2_fill_8 FILLER_0_80_1246 ();
 sg13g2_fill_8 FILLER_0_80_1254 ();
 sg13g2_fill_4 FILLER_0_80_1262 ();
 sg13g2_fill_4 FILLER_0_80_1270 ();
 sg13g2_fill_2 FILLER_0_80_1274 ();
 sg13g2_fill_4 FILLER_0_80_1281 ();
 sg13g2_fill_2 FILLER_0_80_1285 ();
 sg13g2_fill_4 FILLER_0_80_1292 ();
 sg13g2_fill_1 FILLER_0_80_1296 ();
 sg13g2_fill_8 FILLER_0_81_0 ();
 sg13g2_fill_8 FILLER_0_81_8 ();
 sg13g2_fill_8 FILLER_0_81_16 ();
 sg13g2_fill_8 FILLER_0_81_24 ();
 sg13g2_fill_8 FILLER_0_81_32 ();
 sg13g2_fill_8 FILLER_0_81_40 ();
 sg13g2_fill_8 FILLER_0_81_48 ();
 sg13g2_fill_8 FILLER_0_81_56 ();
 sg13g2_fill_8 FILLER_0_81_64 ();
 sg13g2_fill_8 FILLER_0_81_72 ();
 sg13g2_fill_8 FILLER_0_81_80 ();
 sg13g2_fill_8 FILLER_0_81_88 ();
 sg13g2_fill_8 FILLER_0_81_96 ();
 sg13g2_fill_8 FILLER_0_81_104 ();
 sg13g2_fill_8 FILLER_0_81_112 ();
 sg13g2_fill_8 FILLER_0_81_120 ();
 sg13g2_fill_8 FILLER_0_81_128 ();
 sg13g2_fill_8 FILLER_0_81_136 ();
 sg13g2_fill_8 FILLER_0_81_144 ();
 sg13g2_fill_8 FILLER_0_81_152 ();
 sg13g2_fill_8 FILLER_0_81_160 ();
 sg13g2_fill_8 FILLER_0_81_168 ();
 sg13g2_fill_8 FILLER_0_81_176 ();
 sg13g2_fill_8 FILLER_0_81_184 ();
 sg13g2_fill_8 FILLER_0_81_192 ();
 sg13g2_fill_8 FILLER_0_81_200 ();
 sg13g2_fill_8 FILLER_0_81_208 ();
 sg13g2_fill_2 FILLER_0_81_216 ();
 sg13g2_fill_2 FILLER_0_81_223 ();
 sg13g2_fill_8 FILLER_0_81_229 ();
 sg13g2_fill_8 FILLER_0_81_237 ();
 sg13g2_fill_8 FILLER_0_81_245 ();
 sg13g2_fill_8 FILLER_0_81_253 ();
 sg13g2_fill_8 FILLER_0_81_261 ();
 sg13g2_fill_4 FILLER_0_81_269 ();
 sg13g2_fill_8 FILLER_0_81_299 ();
 sg13g2_fill_4 FILLER_0_81_307 ();
 sg13g2_fill_4 FILLER_0_81_337 ();
 sg13g2_fill_1 FILLER_0_81_341 ();
 sg13g2_fill_4 FILLER_0_81_368 ();
 sg13g2_fill_1 FILLER_0_81_372 ();
 sg13g2_fill_4 FILLER_0_81_381 ();
 sg13g2_fill_1 FILLER_0_81_385 ();
 sg13g2_fill_8 FILLER_0_81_391 ();
 sg13g2_fill_2 FILLER_0_81_399 ();
 sg13g2_fill_4 FILLER_0_81_406 ();
 sg13g2_fill_1 FILLER_0_81_410 ();
 sg13g2_fill_2 FILLER_0_81_416 ();
 sg13g2_fill_4 FILLER_0_81_423 ();
 sg13g2_fill_2 FILLER_0_81_432 ();
 sg13g2_fill_4 FILLER_0_81_460 ();
 sg13g2_fill_2 FILLER_0_81_464 ();
 sg13g2_fill_1 FILLER_0_81_466 ();
 sg13g2_fill_2 FILLER_0_81_493 ();
 sg13g2_fill_2 FILLER_0_81_499 ();
 sg13g2_fill_4 FILLER_0_81_511 ();
 sg13g2_fill_2 FILLER_0_81_515 ();
 sg13g2_fill_1 FILLER_0_81_517 ();
 sg13g2_fill_4 FILLER_0_81_524 ();
 sg13g2_fill_2 FILLER_0_81_528 ();
 sg13g2_fill_1 FILLER_0_81_530 ();
 sg13g2_fill_4 FILLER_0_81_535 ();
 sg13g2_fill_1 FILLER_0_81_539 ();
 sg13g2_fill_8 FILLER_0_81_544 ();
 sg13g2_fill_8 FILLER_0_81_552 ();
 sg13g2_fill_4 FILLER_0_81_560 ();
 sg13g2_fill_2 FILLER_0_81_574 ();
 sg13g2_fill_8 FILLER_0_81_581 ();
 sg13g2_fill_1 FILLER_0_81_589 ();
 sg13g2_fill_4 FILLER_0_81_595 ();
 sg13g2_fill_2 FILLER_0_81_599 ();
 sg13g2_fill_8 FILLER_0_81_627 ();
 sg13g2_fill_8 FILLER_0_81_635 ();
 sg13g2_fill_4 FILLER_0_81_643 ();
 sg13g2_fill_4 FILLER_0_81_652 ();
 sg13g2_fill_2 FILLER_0_81_656 ();
 sg13g2_fill_1 FILLER_0_81_658 ();
 sg13g2_fill_2 FILLER_0_81_685 ();
 sg13g2_fill_2 FILLER_0_81_697 ();
 sg13g2_fill_8 FILLER_0_81_704 ();
 sg13g2_fill_1 FILLER_0_81_712 ();
 sg13g2_fill_8 FILLER_0_81_739 ();
 sg13g2_fill_2 FILLER_0_81_752 ();
 sg13g2_fill_2 FILLER_0_81_780 ();
 sg13g2_fill_4 FILLER_0_81_787 ();
 sg13g2_fill_4 FILLER_0_81_801 ();
 sg13g2_fill_2 FILLER_0_81_805 ();
 sg13g2_fill_1 FILLER_0_81_807 ();
 sg13g2_fill_8 FILLER_0_81_813 ();
 sg13g2_fill_2 FILLER_0_81_821 ();
 sg13g2_fill_2 FILLER_0_81_827 ();
 sg13g2_fill_8 FILLER_0_81_834 ();
 sg13g2_fill_8 FILLER_0_81_842 ();
 sg13g2_fill_8 FILLER_0_81_850 ();
 sg13g2_fill_8 FILLER_0_81_858 ();
 sg13g2_fill_8 FILLER_0_81_866 ();
 sg13g2_fill_2 FILLER_0_81_874 ();
 sg13g2_fill_8 FILLER_0_81_882 ();
 sg13g2_fill_2 FILLER_0_81_890 ();
 sg13g2_fill_1 FILLER_0_81_892 ();
 sg13g2_fill_2 FILLER_0_81_903 ();
 sg13g2_fill_8 FILLER_0_81_915 ();
 sg13g2_fill_8 FILLER_0_81_923 ();
 sg13g2_fill_8 FILLER_0_81_931 ();
 sg13g2_fill_8 FILLER_0_81_939 ();
 sg13g2_fill_8 FILLER_0_81_947 ();
 sg13g2_fill_8 FILLER_0_81_955 ();
 sg13g2_fill_8 FILLER_0_81_963 ();
 sg13g2_fill_1 FILLER_0_81_971 ();
 sg13g2_fill_8 FILLER_0_81_977 ();
 sg13g2_fill_8 FILLER_0_81_985 ();
 sg13g2_fill_8 FILLER_0_81_993 ();
 sg13g2_fill_8 FILLER_0_81_1001 ();
 sg13g2_fill_4 FILLER_0_81_1012 ();
 sg13g2_fill_1 FILLER_0_81_1016 ();
 sg13g2_fill_8 FILLER_0_81_1022 ();
 sg13g2_fill_2 FILLER_0_81_1034 ();
 sg13g2_fill_2 FILLER_0_81_1039 ();
 sg13g2_fill_2 FILLER_0_81_1048 ();
 sg13g2_fill_8 FILLER_0_81_1055 ();
 sg13g2_fill_8 FILLER_0_81_1063 ();
 sg13g2_fill_8 FILLER_0_81_1071 ();
 sg13g2_fill_8 FILLER_0_81_1079 ();
 sg13g2_fill_8 FILLER_0_81_1087 ();
 sg13g2_fill_8 FILLER_0_81_1095 ();
 sg13g2_fill_2 FILLER_0_81_1103 ();
 sg13g2_fill_1 FILLER_0_81_1105 ();
 sg13g2_fill_8 FILLER_0_81_1110 ();
 sg13g2_fill_8 FILLER_0_81_1118 ();
 sg13g2_fill_4 FILLER_0_81_1126 ();
 sg13g2_fill_1 FILLER_0_81_1130 ();
 sg13g2_fill_8 FILLER_0_81_1136 ();
 sg13g2_fill_8 FILLER_0_81_1144 ();
 sg13g2_fill_2 FILLER_0_81_1152 ();
 sg13g2_fill_1 FILLER_0_81_1154 ();
 sg13g2_fill_8 FILLER_0_81_1159 ();
 sg13g2_fill_4 FILLER_0_81_1167 ();
 sg13g2_fill_1 FILLER_0_81_1171 ();
 sg13g2_fill_8 FILLER_0_81_1176 ();
 sg13g2_fill_8 FILLER_0_81_1184 ();
 sg13g2_fill_2 FILLER_0_81_1192 ();
 sg13g2_fill_1 FILLER_0_81_1194 ();
 sg13g2_fill_2 FILLER_0_81_1200 ();
 sg13g2_fill_2 FILLER_0_81_1207 ();
 sg13g2_fill_8 FILLER_0_81_1216 ();
 sg13g2_fill_8 FILLER_0_81_1224 ();
 sg13g2_fill_8 FILLER_0_81_1237 ();
 sg13g2_fill_1 FILLER_0_81_1245 ();
 sg13g2_fill_2 FILLER_0_81_1256 ();
 sg13g2_fill_2 FILLER_0_81_1284 ();
 sg13g2_fill_2 FILLER_0_81_1290 ();
 sg13g2_fill_1 FILLER_0_81_1296 ();
 sg13g2_fill_8 FILLER_0_82_0 ();
 sg13g2_fill_8 FILLER_0_82_8 ();
 sg13g2_fill_8 FILLER_0_82_16 ();
 sg13g2_fill_8 FILLER_0_82_24 ();
 sg13g2_fill_8 FILLER_0_82_32 ();
 sg13g2_fill_8 FILLER_0_82_40 ();
 sg13g2_fill_8 FILLER_0_82_48 ();
 sg13g2_fill_8 FILLER_0_82_56 ();
 sg13g2_fill_8 FILLER_0_82_64 ();
 sg13g2_fill_8 FILLER_0_82_72 ();
 sg13g2_fill_8 FILLER_0_82_80 ();
 sg13g2_fill_8 FILLER_0_82_88 ();
 sg13g2_fill_8 FILLER_0_82_96 ();
 sg13g2_fill_8 FILLER_0_82_104 ();
 sg13g2_fill_8 FILLER_0_82_112 ();
 sg13g2_fill_8 FILLER_0_82_120 ();
 sg13g2_fill_8 FILLER_0_82_128 ();
 sg13g2_fill_8 FILLER_0_82_136 ();
 sg13g2_fill_8 FILLER_0_82_144 ();
 sg13g2_fill_8 FILLER_0_82_152 ();
 sg13g2_fill_8 FILLER_0_82_160 ();
 sg13g2_fill_8 FILLER_0_82_168 ();
 sg13g2_fill_8 FILLER_0_82_176 ();
 sg13g2_fill_8 FILLER_0_82_184 ();
 sg13g2_fill_8 FILLER_0_82_192 ();
 sg13g2_fill_8 FILLER_0_82_200 ();
 sg13g2_fill_8 FILLER_0_82_208 ();
 sg13g2_fill_8 FILLER_0_82_216 ();
 sg13g2_fill_8 FILLER_0_82_224 ();
 sg13g2_fill_8 FILLER_0_82_232 ();
 sg13g2_fill_8 FILLER_0_82_240 ();
 sg13g2_fill_8 FILLER_0_82_248 ();
 sg13g2_fill_2 FILLER_0_82_256 ();
 sg13g2_fill_1 FILLER_0_82_258 ();
 sg13g2_fill_8 FILLER_0_82_285 ();
 sg13g2_fill_8 FILLER_0_82_293 ();
 sg13g2_fill_8 FILLER_0_82_305 ();
 sg13g2_fill_8 FILLER_0_82_318 ();
 sg13g2_fill_4 FILLER_0_82_330 ();
 sg13g2_fill_2 FILLER_0_82_339 ();
 sg13g2_fill_8 FILLER_0_82_362 ();
 sg13g2_fill_8 FILLER_0_82_370 ();
 sg13g2_fill_4 FILLER_0_82_378 ();
 sg13g2_fill_2 FILLER_0_82_382 ();
 sg13g2_fill_8 FILLER_0_82_389 ();
 sg13g2_fill_8 FILLER_0_82_397 ();
 sg13g2_fill_8 FILLER_0_82_405 ();
 sg13g2_fill_2 FILLER_0_82_418 ();
 sg13g2_fill_2 FILLER_0_82_425 ();
 sg13g2_fill_8 FILLER_0_82_432 ();
 sg13g2_fill_8 FILLER_0_82_440 ();
 sg13g2_fill_8 FILLER_0_82_448 ();
 sg13g2_fill_4 FILLER_0_82_456 ();
 sg13g2_fill_4 FILLER_0_82_465 ();
 sg13g2_fill_2 FILLER_0_82_474 ();
 sg13g2_fill_2 FILLER_0_82_502 ();
 sg13g2_fill_1 FILLER_0_82_504 ();
 sg13g2_fill_2 FILLER_0_82_515 ();
 sg13g2_fill_1 FILLER_0_82_517 ();
 sg13g2_fill_4 FILLER_0_82_522 ();
 sg13g2_fill_2 FILLER_0_82_530 ();
 sg13g2_fill_2 FILLER_0_82_537 ();
 sg13g2_fill_4 FILLER_0_82_565 ();
 sg13g2_fill_1 FILLER_0_82_569 ();
 sg13g2_fill_2 FILLER_0_82_574 ();
 sg13g2_fill_8 FILLER_0_82_582 ();
 sg13g2_fill_8 FILLER_0_82_590 ();
 sg13g2_fill_4 FILLER_0_82_604 ();
 sg13g2_fill_2 FILLER_0_82_608 ();
 sg13g2_fill_1 FILLER_0_82_610 ();
 sg13g2_fill_2 FILLER_0_82_615 ();
 sg13g2_fill_4 FILLER_0_82_643 ();
 sg13g2_fill_2 FILLER_0_82_647 ();
 sg13g2_fill_8 FILLER_0_82_654 ();
 sg13g2_fill_8 FILLER_0_82_662 ();
 sg13g2_fill_8 FILLER_0_82_670 ();
 sg13g2_fill_8 FILLER_0_82_678 ();
 sg13g2_fill_4 FILLER_0_82_686 ();
 sg13g2_fill_4 FILLER_0_82_700 ();
 sg13g2_fill_2 FILLER_0_82_704 ();
 sg13g2_fill_1 FILLER_0_82_706 ();
 sg13g2_fill_8 FILLER_0_82_713 ();
 sg13g2_fill_8 FILLER_0_82_721 ();
 sg13g2_fill_1 FILLER_0_82_729 ();
 sg13g2_fill_8 FILLER_0_82_734 ();
 sg13g2_fill_2 FILLER_0_82_742 ();
 sg13g2_fill_2 FILLER_0_82_749 ();
 sg13g2_fill_2 FILLER_0_82_756 ();
 sg13g2_fill_2 FILLER_0_82_763 ();
 sg13g2_fill_4 FILLER_0_82_770 ();
 sg13g2_fill_1 FILLER_0_82_774 ();
 sg13g2_fill_4 FILLER_0_82_780 ();
 sg13g2_fill_2 FILLER_0_82_790 ();
 sg13g2_fill_1 FILLER_0_82_792 ();
 sg13g2_fill_2 FILLER_0_82_819 ();
 sg13g2_fill_2 FILLER_0_82_826 ();
 sg13g2_fill_2 FILLER_0_82_834 ();
 sg13g2_fill_4 FILLER_0_82_842 ();
 sg13g2_fill_2 FILLER_0_82_846 ();
 sg13g2_fill_2 FILLER_0_82_857 ();
 sg13g2_fill_4 FILLER_0_82_865 ();
 sg13g2_fill_2 FILLER_0_82_869 ();
 sg13g2_fill_8 FILLER_0_82_876 ();
 sg13g2_fill_2 FILLER_0_82_884 ();
 sg13g2_fill_1 FILLER_0_82_886 ();
 sg13g2_fill_2 FILLER_0_82_897 ();
 sg13g2_fill_4 FILLER_0_82_909 ();
 sg13g2_fill_2 FILLER_0_82_917 ();
 sg13g2_fill_1 FILLER_0_82_919 ();
 sg13g2_fill_2 FILLER_0_82_925 ();
 sg13g2_fill_4 FILLER_0_82_933 ();
 sg13g2_fill_2 FILLER_0_82_937 ();
 sg13g2_fill_1 FILLER_0_82_939 ();
 sg13g2_fill_8 FILLER_0_82_944 ();
 sg13g2_fill_8 FILLER_0_82_952 ();
 sg13g2_fill_8 FILLER_0_82_960 ();
 sg13g2_fill_4 FILLER_0_82_968 ();
 sg13g2_fill_2 FILLER_0_82_977 ();
 sg13g2_fill_2 FILLER_0_82_985 ();
 sg13g2_fill_4 FILLER_0_82_992 ();
 sg13g2_fill_1 FILLER_0_82_996 ();
 sg13g2_fill_4 FILLER_0_82_1003 ();
 sg13g2_fill_2 FILLER_0_82_1007 ();
 sg13g2_fill_4 FILLER_0_82_1015 ();
 sg13g2_fill_2 FILLER_0_82_1019 ();
 sg13g2_fill_8 FILLER_0_82_1026 ();
 sg13g2_fill_8 FILLER_0_82_1034 ();
 sg13g2_fill_4 FILLER_0_82_1042 ();
 sg13g2_fill_4 FILLER_0_82_1051 ();
 sg13g2_fill_2 FILLER_0_82_1055 ();
 sg13g2_fill_1 FILLER_0_82_1057 ();
 sg13g2_fill_8 FILLER_0_82_1062 ();
 sg13g2_fill_8 FILLER_0_82_1070 ();
 sg13g2_fill_4 FILLER_0_82_1078 ();
 sg13g2_fill_1 FILLER_0_82_1082 ();
 sg13g2_fill_2 FILLER_0_82_1086 ();
 sg13g2_fill_8 FILLER_0_82_1093 ();
 sg13g2_fill_8 FILLER_0_82_1101 ();
 sg13g2_fill_8 FILLER_0_82_1109 ();
 sg13g2_fill_8 FILLER_0_82_1117 ();
 sg13g2_fill_8 FILLER_0_82_1125 ();
 sg13g2_fill_8 FILLER_0_82_1133 ();
 sg13g2_fill_2 FILLER_0_82_1141 ();
 sg13g2_fill_2 FILLER_0_82_1147 ();
 sg13g2_fill_2 FILLER_0_82_1153 ();
 sg13g2_fill_2 FILLER_0_82_1160 ();
 sg13g2_fill_1 FILLER_0_82_1162 ();
 sg13g2_fill_2 FILLER_0_82_1170 ();
 sg13g2_fill_8 FILLER_0_82_1177 ();
 sg13g2_fill_2 FILLER_0_82_1185 ();
 sg13g2_fill_1 FILLER_0_82_1187 ();
 sg13g2_fill_8 FILLER_0_82_1193 ();
 sg13g2_fill_4 FILLER_0_82_1201 ();
 sg13g2_fill_2 FILLER_0_82_1205 ();
 sg13g2_fill_2 FILLER_0_82_1214 ();
 sg13g2_fill_8 FILLER_0_82_1221 ();
 sg13g2_fill_2 FILLER_0_82_1229 ();
 sg13g2_fill_1 FILLER_0_82_1231 ();
 sg13g2_fill_4 FILLER_0_82_1236 ();
 sg13g2_fill_1 FILLER_0_82_1240 ();
 sg13g2_fill_2 FILLER_0_82_1251 ();
 sg13g2_fill_1 FILLER_0_82_1253 ();
 sg13g2_fill_8 FILLER_0_82_1259 ();
 sg13g2_fill_2 FILLER_0_82_1267 ();
 sg13g2_fill_2 FILLER_0_82_1274 ();
 sg13g2_fill_2 FILLER_0_82_1284 ();
 sg13g2_fill_2 FILLER_0_82_1290 ();
 sg13g2_fill_1 FILLER_0_82_1296 ();
 sg13g2_fill_8 FILLER_0_83_0 ();
 sg13g2_fill_8 FILLER_0_83_8 ();
 sg13g2_fill_8 FILLER_0_83_16 ();
 sg13g2_fill_8 FILLER_0_83_24 ();
 sg13g2_fill_8 FILLER_0_83_32 ();
 sg13g2_fill_8 FILLER_0_83_40 ();
 sg13g2_fill_8 FILLER_0_83_48 ();
 sg13g2_fill_8 FILLER_0_83_56 ();
 sg13g2_fill_8 FILLER_0_83_64 ();
 sg13g2_fill_8 FILLER_0_83_72 ();
 sg13g2_fill_8 FILLER_0_83_80 ();
 sg13g2_fill_8 FILLER_0_83_88 ();
 sg13g2_fill_8 FILLER_0_83_96 ();
 sg13g2_fill_8 FILLER_0_83_104 ();
 sg13g2_fill_8 FILLER_0_83_112 ();
 sg13g2_fill_8 FILLER_0_83_120 ();
 sg13g2_fill_8 FILLER_0_83_128 ();
 sg13g2_fill_8 FILLER_0_83_136 ();
 sg13g2_fill_8 FILLER_0_83_144 ();
 sg13g2_fill_8 FILLER_0_83_152 ();
 sg13g2_fill_8 FILLER_0_83_160 ();
 sg13g2_fill_8 FILLER_0_83_168 ();
 sg13g2_fill_8 FILLER_0_83_176 ();
 sg13g2_fill_8 FILLER_0_83_184 ();
 sg13g2_fill_8 FILLER_0_83_192 ();
 sg13g2_fill_8 FILLER_0_83_200 ();
 sg13g2_fill_8 FILLER_0_83_208 ();
 sg13g2_fill_8 FILLER_0_83_216 ();
 sg13g2_fill_8 FILLER_0_83_224 ();
 sg13g2_fill_8 FILLER_0_83_232 ();
 sg13g2_fill_8 FILLER_0_83_240 ();
 sg13g2_fill_8 FILLER_0_83_248 ();
 sg13g2_fill_8 FILLER_0_83_256 ();
 sg13g2_fill_8 FILLER_0_83_264 ();
 sg13g2_fill_2 FILLER_0_83_277 ();
 sg13g2_fill_2 FILLER_0_83_283 ();
 sg13g2_fill_1 FILLER_0_83_285 ();
 sg13g2_fill_8 FILLER_0_83_292 ();
 sg13g2_fill_4 FILLER_0_83_300 ();
 sg13g2_fill_2 FILLER_0_83_304 ();
 sg13g2_fill_4 FILLER_0_83_311 ();
 sg13g2_fill_1 FILLER_0_83_315 ();
 sg13g2_fill_2 FILLER_0_83_321 ();
 sg13g2_fill_2 FILLER_0_83_349 ();
 sg13g2_fill_8 FILLER_0_83_355 ();
 sg13g2_fill_8 FILLER_0_83_363 ();
 sg13g2_fill_8 FILLER_0_83_371 ();
 sg13g2_fill_4 FILLER_0_83_379 ();
 sg13g2_fill_1 FILLER_0_83_383 ();
 sg13g2_fill_2 FILLER_0_83_389 ();
 sg13g2_fill_8 FILLER_0_83_395 ();
 sg13g2_fill_8 FILLER_0_83_429 ();
 sg13g2_fill_8 FILLER_0_83_437 ();
 sg13g2_fill_8 FILLER_0_83_445 ();
 sg13g2_fill_8 FILLER_0_83_453 ();
 sg13g2_fill_8 FILLER_0_83_461 ();
 sg13g2_fill_4 FILLER_0_83_469 ();
 sg13g2_fill_2 FILLER_0_83_477 ();
 sg13g2_fill_4 FILLER_0_83_484 ();
 sg13g2_fill_2 FILLER_0_83_488 ();
 sg13g2_fill_1 FILLER_0_83_490 ();
 sg13g2_fill_8 FILLER_0_83_496 ();
 sg13g2_fill_8 FILLER_0_83_504 ();
 sg13g2_fill_8 FILLER_0_83_512 ();
 sg13g2_fill_8 FILLER_0_83_520 ();
 sg13g2_fill_8 FILLER_0_83_528 ();
 sg13g2_fill_8 FILLER_0_83_536 ();
 sg13g2_fill_4 FILLER_0_83_544 ();
 sg13g2_fill_8 FILLER_0_83_553 ();
 sg13g2_fill_8 FILLER_0_83_561 ();
 sg13g2_fill_2 FILLER_0_83_569 ();
 sg13g2_fill_1 FILLER_0_83_571 ();
 sg13g2_fill_2 FILLER_0_83_576 ();
 sg13g2_fill_8 FILLER_0_83_583 ();
 sg13g2_fill_4 FILLER_0_83_591 ();
 sg13g2_fill_2 FILLER_0_83_595 ();
 sg13g2_fill_2 FILLER_0_83_603 ();
 sg13g2_fill_2 FILLER_0_83_611 ();
 sg13g2_fill_2 FILLER_0_83_617 ();
 sg13g2_fill_1 FILLER_0_83_619 ();
 sg13g2_fill_4 FILLER_0_83_626 ();
 sg13g2_fill_2 FILLER_0_83_635 ();
 sg13g2_fill_8 FILLER_0_83_642 ();
 sg13g2_fill_8 FILLER_0_83_654 ();
 sg13g2_fill_1 FILLER_0_83_662 ();
 sg13g2_fill_2 FILLER_0_83_668 ();
 sg13g2_fill_1 FILLER_0_83_670 ();
 sg13g2_fill_2 FILLER_0_83_697 ();
 sg13g2_fill_8 FILLER_0_83_703 ();
 sg13g2_fill_4 FILLER_0_83_711 ();
 sg13g2_fill_8 FILLER_0_83_719 ();
 sg13g2_fill_8 FILLER_0_83_727 ();
 sg13g2_fill_2 FILLER_0_83_735 ();
 sg13g2_fill_8 FILLER_0_83_742 ();
 sg13g2_fill_2 FILLER_0_83_776 ();
 sg13g2_fill_8 FILLER_0_83_788 ();
 sg13g2_fill_4 FILLER_0_83_800 ();
 sg13g2_fill_2 FILLER_0_83_809 ();
 sg13g2_fill_2 FILLER_0_83_816 ();
 sg13g2_fill_1 FILLER_0_83_818 ();
 sg13g2_fill_8 FILLER_0_83_825 ();
 sg13g2_fill_1 FILLER_0_83_833 ();
 sg13g2_fill_8 FILLER_0_83_838 ();
 sg13g2_fill_8 FILLER_0_83_850 ();
 sg13g2_fill_8 FILLER_0_83_858 ();
 sg13g2_fill_8 FILLER_0_83_866 ();
 sg13g2_fill_4 FILLER_0_83_874 ();
 sg13g2_fill_2 FILLER_0_83_878 ();
 sg13g2_fill_1 FILLER_0_83_880 ();
 sg13g2_fill_8 FILLER_0_83_886 ();
 sg13g2_fill_4 FILLER_0_83_894 ();
 sg13g2_fill_4 FILLER_0_83_908 ();
 sg13g2_fill_1 FILLER_0_83_912 ();
 sg13g2_fill_8 FILLER_0_83_918 ();
 sg13g2_fill_2 FILLER_0_83_926 ();
 sg13g2_fill_1 FILLER_0_83_928 ();
 sg13g2_fill_2 FILLER_0_83_933 ();
 sg13g2_fill_4 FILLER_0_83_939 ();
 sg13g2_fill_2 FILLER_0_83_943 ();
 sg13g2_fill_1 FILLER_0_83_945 ();
 sg13g2_fill_4 FILLER_0_83_951 ();
 sg13g2_fill_1 FILLER_0_83_955 ();
 sg13g2_fill_2 FILLER_0_83_964 ();
 sg13g2_fill_8 FILLER_0_83_972 ();
 sg13g2_fill_4 FILLER_0_83_984 ();
 sg13g2_fill_1 FILLER_0_83_988 ();
 sg13g2_fill_2 FILLER_0_83_994 ();
 sg13g2_fill_4 FILLER_0_83_1001 ();
 sg13g2_fill_1 FILLER_0_83_1005 ();
 sg13g2_fill_2 FILLER_0_83_1011 ();
 sg13g2_fill_1 FILLER_0_83_1013 ();
 sg13g2_fill_8 FILLER_0_83_1019 ();
 sg13g2_fill_4 FILLER_0_83_1027 ();
 sg13g2_fill_2 FILLER_0_83_1037 ();
 sg13g2_fill_2 FILLER_0_83_1043 ();
 sg13g2_fill_4 FILLER_0_83_1051 ();
 sg13g2_fill_2 FILLER_0_83_1059 ();
 sg13g2_fill_4 FILLER_0_83_1067 ();
 sg13g2_fill_1 FILLER_0_83_1071 ();
 sg13g2_fill_4 FILLER_0_83_1077 ();
 sg13g2_fill_4 FILLER_0_83_1086 ();
 sg13g2_fill_1 FILLER_0_83_1090 ();
 sg13g2_fill_8 FILLER_0_83_1096 ();
 sg13g2_fill_2 FILLER_0_83_1104 ();
 sg13g2_fill_2 FILLER_0_83_1111 ();
 sg13g2_fill_2 FILLER_0_83_1116 ();
 sg13g2_fill_8 FILLER_0_83_1124 ();
 sg13g2_fill_2 FILLER_0_83_1132 ();
 sg13g2_fill_8 FILLER_0_83_1138 ();
 sg13g2_fill_2 FILLER_0_83_1151 ();
 sg13g2_fill_1 FILLER_0_83_1153 ();
 sg13g2_fill_2 FILLER_0_83_1161 ();
 sg13g2_fill_1 FILLER_0_83_1163 ();
 sg13g2_fill_2 FILLER_0_83_1169 ();
 sg13g2_fill_1 FILLER_0_83_1171 ();
 sg13g2_fill_2 FILLER_0_83_1180 ();
 sg13g2_fill_1 FILLER_0_83_1182 ();
 sg13g2_fill_4 FILLER_0_83_1190 ();
 sg13g2_fill_2 FILLER_0_83_1200 ();
 sg13g2_fill_2 FILLER_0_83_1206 ();
 sg13g2_fill_2 FILLER_0_83_1212 ();
 sg13g2_fill_2 FILLER_0_83_1218 ();
 sg13g2_fill_8 FILLER_0_83_1224 ();
 sg13g2_fill_2 FILLER_0_83_1236 ();
 sg13g2_fill_2 FILLER_0_83_1243 ();
 sg13g2_fill_4 FILLER_0_83_1251 ();
 sg13g2_fill_2 FILLER_0_83_1255 ();
 sg13g2_fill_4 FILLER_0_83_1262 ();
 sg13g2_fill_2 FILLER_0_83_1271 ();
 sg13g2_fill_8 FILLER_0_83_1278 ();
 sg13g2_fill_4 FILLER_0_83_1286 ();
 sg13g2_fill_2 FILLER_0_83_1290 ();
 sg13g2_fill_1 FILLER_0_83_1296 ();
 sg13g2_fill_8 FILLER_0_84_0 ();
 sg13g2_fill_8 FILLER_0_84_8 ();
 sg13g2_fill_8 FILLER_0_84_16 ();
 sg13g2_fill_8 FILLER_0_84_24 ();
 sg13g2_fill_8 FILLER_0_84_32 ();
 sg13g2_fill_8 FILLER_0_84_40 ();
 sg13g2_fill_8 FILLER_0_84_48 ();
 sg13g2_fill_8 FILLER_0_84_56 ();
 sg13g2_fill_8 FILLER_0_84_64 ();
 sg13g2_fill_8 FILLER_0_84_72 ();
 sg13g2_fill_8 FILLER_0_84_80 ();
 sg13g2_fill_8 FILLER_0_84_88 ();
 sg13g2_fill_8 FILLER_0_84_96 ();
 sg13g2_fill_8 FILLER_0_84_104 ();
 sg13g2_fill_8 FILLER_0_84_112 ();
 sg13g2_fill_8 FILLER_0_84_120 ();
 sg13g2_fill_8 FILLER_0_84_128 ();
 sg13g2_fill_8 FILLER_0_84_136 ();
 sg13g2_fill_8 FILLER_0_84_144 ();
 sg13g2_fill_8 FILLER_0_84_152 ();
 sg13g2_fill_8 FILLER_0_84_160 ();
 sg13g2_fill_8 FILLER_0_84_168 ();
 sg13g2_fill_8 FILLER_0_84_176 ();
 sg13g2_fill_8 FILLER_0_84_184 ();
 sg13g2_fill_8 FILLER_0_84_192 ();
 sg13g2_fill_8 FILLER_0_84_200 ();
 sg13g2_fill_8 FILLER_0_84_208 ();
 sg13g2_fill_8 FILLER_0_84_216 ();
 sg13g2_fill_4 FILLER_0_84_224 ();
 sg13g2_fill_2 FILLER_0_84_233 ();
 sg13g2_fill_2 FILLER_0_84_239 ();
 sg13g2_fill_4 FILLER_0_84_246 ();
 sg13g2_fill_2 FILLER_0_84_250 ();
 sg13g2_fill_2 FILLER_0_84_257 ();
 sg13g2_fill_8 FILLER_0_84_266 ();
 sg13g2_fill_8 FILLER_0_84_274 ();
 sg13g2_fill_8 FILLER_0_84_282 ();
 sg13g2_fill_4 FILLER_0_84_290 ();
 sg13g2_fill_8 FILLER_0_84_299 ();
 sg13g2_fill_4 FILLER_0_84_307 ();
 sg13g2_fill_8 FILLER_0_84_319 ();
 sg13g2_fill_8 FILLER_0_84_327 ();
 sg13g2_fill_8 FILLER_0_84_335 ();
 sg13g2_fill_2 FILLER_0_84_343 ();
 sg13g2_fill_1 FILLER_0_84_345 ();
 sg13g2_fill_8 FILLER_0_84_351 ();
 sg13g2_fill_4 FILLER_0_84_359 ();
 sg13g2_fill_1 FILLER_0_84_363 ();
 sg13g2_fill_2 FILLER_0_84_371 ();
 sg13g2_fill_2 FILLER_0_84_399 ();
 sg13g2_fill_2 FILLER_0_84_406 ();
 sg13g2_fill_1 FILLER_0_84_408 ();
 sg13g2_fill_2 FILLER_0_84_413 ();
 sg13g2_fill_1 FILLER_0_84_415 ();
 sg13g2_fill_4 FILLER_0_84_421 ();
 sg13g2_fill_4 FILLER_0_84_429 ();
 sg13g2_fill_2 FILLER_0_84_433 ();
 sg13g2_fill_8 FILLER_0_84_442 ();
 sg13g2_fill_8 FILLER_0_84_450 ();
 sg13g2_fill_8 FILLER_0_84_458 ();
 sg13g2_fill_8 FILLER_0_84_472 ();
 sg13g2_fill_8 FILLER_0_84_480 ();
 sg13g2_fill_8 FILLER_0_84_488 ();
 sg13g2_fill_8 FILLER_0_84_496 ();
 sg13g2_fill_8 FILLER_0_84_504 ();
 sg13g2_fill_8 FILLER_0_84_512 ();
 sg13g2_fill_8 FILLER_0_84_520 ();
 sg13g2_fill_4 FILLER_0_84_528 ();
 sg13g2_fill_1 FILLER_0_84_532 ();
 sg13g2_fill_8 FILLER_0_84_537 ();
 sg13g2_fill_8 FILLER_0_84_545 ();
 sg13g2_fill_8 FILLER_0_84_553 ();
 sg13g2_fill_4 FILLER_0_84_561 ();
 sg13g2_fill_2 FILLER_0_84_565 ();
 sg13g2_fill_1 FILLER_0_84_567 ();
 sg13g2_fill_8 FILLER_0_84_574 ();
 sg13g2_fill_8 FILLER_0_84_582 ();
 sg13g2_fill_8 FILLER_0_84_590 ();
 sg13g2_fill_8 FILLER_0_84_598 ();
 sg13g2_fill_1 FILLER_0_84_606 ();
 sg13g2_fill_8 FILLER_0_84_612 ();
 sg13g2_fill_8 FILLER_0_84_620 ();
 sg13g2_fill_8 FILLER_0_84_628 ();
 sg13g2_fill_8 FILLER_0_84_636 ();
 sg13g2_fill_8 FILLER_0_84_644 ();
 sg13g2_fill_8 FILLER_0_84_652 ();
 sg13g2_fill_8 FILLER_0_84_670 ();
 sg13g2_fill_1 FILLER_0_84_678 ();
 sg13g2_fill_2 FILLER_0_84_700 ();
 sg13g2_fill_8 FILLER_0_84_708 ();
 sg13g2_fill_2 FILLER_0_84_716 ();
 sg13g2_fill_4 FILLER_0_84_723 ();
 sg13g2_fill_1 FILLER_0_84_727 ();
 sg13g2_fill_2 FILLER_0_84_733 ();
 sg13g2_fill_2 FILLER_0_84_761 ();
 sg13g2_fill_8 FILLER_0_84_768 ();
 sg13g2_fill_8 FILLER_0_84_776 ();
 sg13g2_fill_1 FILLER_0_84_784 ();
 sg13g2_fill_2 FILLER_0_84_795 ();
 sg13g2_fill_4 FILLER_0_84_823 ();
 sg13g2_fill_2 FILLER_0_84_833 ();
 sg13g2_fill_1 FILLER_0_84_835 ();
 sg13g2_fill_4 FILLER_0_84_841 ();
 sg13g2_fill_2 FILLER_0_84_845 ();
 sg13g2_fill_2 FILLER_0_84_851 ();
 sg13g2_fill_1 FILLER_0_84_853 ();
 sg13g2_fill_2 FILLER_0_84_858 ();
 sg13g2_fill_2 FILLER_0_84_866 ();
 sg13g2_fill_8 FILLER_0_84_873 ();
 sg13g2_fill_8 FILLER_0_84_881 ();
 sg13g2_fill_8 FILLER_0_84_889 ();
 sg13g2_fill_8 FILLER_0_84_907 ();
 sg13g2_fill_1 FILLER_0_84_915 ();
 sg13g2_fill_8 FILLER_0_84_926 ();
 sg13g2_fill_8 FILLER_0_84_934 ();
 sg13g2_fill_2 FILLER_0_84_942 ();
 sg13g2_fill_8 FILLER_0_84_950 ();
 sg13g2_fill_8 FILLER_0_84_958 ();
 sg13g2_fill_8 FILLER_0_84_966 ();
 sg13g2_fill_1 FILLER_0_84_974 ();
 sg13g2_fill_4 FILLER_0_84_979 ();
 sg13g2_fill_1 FILLER_0_84_983 ();
 sg13g2_fill_2 FILLER_0_84_989 ();
 sg13g2_fill_1 FILLER_0_84_991 ();
 sg13g2_fill_2 FILLER_0_84_996 ();
 sg13g2_fill_2 FILLER_0_84_1003 ();
 sg13g2_fill_2 FILLER_0_84_1010 ();
 sg13g2_fill_2 FILLER_0_84_1017 ();
 sg13g2_fill_2 FILLER_0_84_1023 ();
 sg13g2_fill_2 FILLER_0_84_1030 ();
 sg13g2_fill_4 FILLER_0_84_1036 ();
 sg13g2_fill_2 FILLER_0_84_1045 ();
 sg13g2_fill_2 FILLER_0_84_1054 ();
 sg13g2_fill_2 FILLER_0_84_1061 ();
 sg13g2_fill_2 FILLER_0_84_1067 ();
 sg13g2_fill_1 FILLER_0_84_1069 ();
 sg13g2_fill_4 FILLER_0_84_1074 ();
 sg13g2_fill_1 FILLER_0_84_1078 ();
 sg13g2_fill_2 FILLER_0_84_1086 ();
 sg13g2_fill_4 FILLER_0_84_1096 ();
 sg13g2_fill_1 FILLER_0_84_1100 ();
 sg13g2_fill_8 FILLER_0_84_1106 ();
 sg13g2_fill_8 FILLER_0_84_1114 ();
 sg13g2_fill_4 FILLER_0_84_1126 ();
 sg13g2_fill_2 FILLER_0_84_1135 ();
 sg13g2_fill_2 FILLER_0_84_1142 ();
 sg13g2_fill_4 FILLER_0_84_1149 ();
 sg13g2_fill_4 FILLER_0_84_1158 ();
 sg13g2_fill_2 FILLER_0_84_1166 ();
 sg13g2_fill_1 FILLER_0_84_1168 ();
 sg13g2_fill_2 FILLER_0_84_1174 ();
 sg13g2_fill_4 FILLER_0_84_1181 ();
 sg13g2_fill_2 FILLER_0_84_1185 ();
 sg13g2_fill_2 FILLER_0_84_1192 ();
 sg13g2_fill_2 FILLER_0_84_1201 ();
 sg13g2_fill_2 FILLER_0_84_1208 ();
 sg13g2_fill_4 FILLER_0_84_1215 ();
 sg13g2_fill_2 FILLER_0_84_1219 ();
 sg13g2_fill_1 FILLER_0_84_1221 ();
 sg13g2_fill_4 FILLER_0_84_1227 ();
 sg13g2_fill_2 FILLER_0_84_1231 ();
 sg13g2_fill_1 FILLER_0_84_1233 ();
 sg13g2_fill_2 FILLER_0_84_1239 ();
 sg13g2_fill_2 FILLER_0_84_1247 ();
 sg13g2_fill_2 FILLER_0_84_1254 ();
 sg13g2_fill_2 FILLER_0_84_1260 ();
 sg13g2_fill_1 FILLER_0_84_1262 ();
 sg13g2_fill_4 FILLER_0_84_1267 ();
 sg13g2_fill_2 FILLER_0_84_1271 ();
 sg13g2_fill_2 FILLER_0_84_1278 ();
 sg13g2_fill_8 FILLER_0_84_1285 ();
 sg13g2_fill_4 FILLER_0_84_1293 ();
 sg13g2_fill_8 FILLER_0_85_0 ();
 sg13g2_fill_8 FILLER_0_85_8 ();
 sg13g2_fill_8 FILLER_0_85_16 ();
 sg13g2_fill_8 FILLER_0_85_24 ();
 sg13g2_fill_8 FILLER_0_85_32 ();
 sg13g2_fill_8 FILLER_0_85_40 ();
 sg13g2_fill_8 FILLER_0_85_48 ();
 sg13g2_fill_8 FILLER_0_85_56 ();
 sg13g2_fill_8 FILLER_0_85_64 ();
 sg13g2_fill_8 FILLER_0_85_72 ();
 sg13g2_fill_8 FILLER_0_85_80 ();
 sg13g2_fill_8 FILLER_0_85_88 ();
 sg13g2_fill_8 FILLER_0_85_96 ();
 sg13g2_fill_8 FILLER_0_85_104 ();
 sg13g2_fill_8 FILLER_0_85_112 ();
 sg13g2_fill_8 FILLER_0_85_120 ();
 sg13g2_fill_8 FILLER_0_85_128 ();
 sg13g2_fill_8 FILLER_0_85_136 ();
 sg13g2_fill_8 FILLER_0_85_144 ();
 sg13g2_fill_8 FILLER_0_85_152 ();
 sg13g2_fill_8 FILLER_0_85_160 ();
 sg13g2_fill_8 FILLER_0_85_168 ();
 sg13g2_fill_8 FILLER_0_85_176 ();
 sg13g2_fill_8 FILLER_0_85_184 ();
 sg13g2_fill_8 FILLER_0_85_192 ();
 sg13g2_fill_8 FILLER_0_85_200 ();
 sg13g2_fill_4 FILLER_0_85_208 ();
 sg13g2_fill_2 FILLER_0_85_212 ();
 sg13g2_fill_4 FILLER_0_85_240 ();
 sg13g2_fill_8 FILLER_0_85_250 ();
 sg13g2_fill_4 FILLER_0_85_258 ();
 sg13g2_fill_2 FILLER_0_85_262 ();
 sg13g2_fill_1 FILLER_0_85_264 ();
 sg13g2_fill_4 FILLER_0_85_272 ();
 sg13g2_fill_8 FILLER_0_85_282 ();
 sg13g2_fill_8 FILLER_0_85_290 ();
 sg13g2_fill_2 FILLER_0_85_303 ();
 sg13g2_fill_1 FILLER_0_85_305 ();
 sg13g2_fill_4 FILLER_0_85_316 ();
 sg13g2_fill_2 FILLER_0_85_320 ();
 sg13g2_fill_2 FILLER_0_85_327 ();
 sg13g2_fill_1 FILLER_0_85_329 ();
 sg13g2_fill_8 FILLER_0_85_336 ();
 sg13g2_fill_8 FILLER_0_85_344 ();
 sg13g2_fill_8 FILLER_0_85_352 ();
 sg13g2_fill_8 FILLER_0_85_372 ();
 sg13g2_fill_8 FILLER_0_85_380 ();
 sg13g2_fill_8 FILLER_0_85_388 ();
 sg13g2_fill_2 FILLER_0_85_396 ();
 sg13g2_fill_1 FILLER_0_85_398 ();
 sg13g2_fill_2 FILLER_0_85_405 ();
 sg13g2_fill_1 FILLER_0_85_407 ();
 sg13g2_fill_2 FILLER_0_85_414 ();
 sg13g2_fill_2 FILLER_0_85_422 ();
 sg13g2_fill_2 FILLER_0_85_429 ();
 sg13g2_fill_8 FILLER_0_85_438 ();
 sg13g2_fill_8 FILLER_0_85_446 ();
 sg13g2_fill_8 FILLER_0_85_454 ();
 sg13g2_fill_8 FILLER_0_85_462 ();
 sg13g2_fill_8 FILLER_0_85_470 ();
 sg13g2_fill_8 FILLER_0_85_478 ();
 sg13g2_fill_8 FILLER_0_85_486 ();
 sg13g2_fill_8 FILLER_0_85_494 ();
 sg13g2_fill_8 FILLER_0_85_502 ();
 sg13g2_fill_2 FILLER_0_85_510 ();
 sg13g2_fill_2 FILLER_0_85_517 ();
 sg13g2_fill_2 FILLER_0_85_545 ();
 sg13g2_fill_2 FILLER_0_85_552 ();
 sg13g2_fill_4 FILLER_0_85_559 ();
 sg13g2_fill_2 FILLER_0_85_563 ();
 sg13g2_fill_2 FILLER_0_85_570 ();
 sg13g2_fill_8 FILLER_0_85_577 ();
 sg13g2_fill_4 FILLER_0_85_585 ();
 sg13g2_fill_2 FILLER_0_85_589 ();
 sg13g2_fill_8 FILLER_0_85_617 ();
 sg13g2_fill_8 FILLER_0_85_625 ();
 sg13g2_fill_8 FILLER_0_85_633 ();
 sg13g2_fill_2 FILLER_0_85_641 ();
 sg13g2_fill_1 FILLER_0_85_643 ();
 sg13g2_fill_2 FILLER_0_85_654 ();
 sg13g2_fill_8 FILLER_0_85_682 ();
 sg13g2_fill_8 FILLER_0_85_690 ();
 sg13g2_fill_8 FILLER_0_85_698 ();
 sg13g2_fill_4 FILLER_0_85_706 ();
 sg13g2_fill_2 FILLER_0_85_710 ();
 sg13g2_fill_1 FILLER_0_85_712 ();
 sg13g2_fill_8 FILLER_0_85_718 ();
 sg13g2_fill_4 FILLER_0_85_726 ();
 sg13g2_fill_1 FILLER_0_85_730 ();
 sg13g2_fill_4 FILLER_0_85_741 ();
 sg13g2_fill_2 FILLER_0_85_745 ();
 sg13g2_fill_1 FILLER_0_85_747 ();
 sg13g2_fill_2 FILLER_0_85_753 ();
 sg13g2_fill_1 FILLER_0_85_755 ();
 sg13g2_fill_2 FILLER_0_85_761 ();
 sg13g2_fill_8 FILLER_0_85_768 ();
 sg13g2_fill_2 FILLER_0_85_776 ();
 sg13g2_fill_1 FILLER_0_85_778 ();
 sg13g2_fill_2 FILLER_0_85_784 ();
 sg13g2_fill_4 FILLER_0_85_792 ();
 sg13g2_fill_8 FILLER_0_85_801 ();
 sg13g2_fill_8 FILLER_0_85_809 ();
 sg13g2_fill_4 FILLER_0_85_817 ();
 sg13g2_fill_2 FILLER_0_85_821 ();
 sg13g2_fill_1 FILLER_0_85_823 ();
 sg13g2_fill_2 FILLER_0_85_828 ();
 sg13g2_fill_1 FILLER_0_85_830 ();
 sg13g2_fill_2 FILLER_0_85_835 ();
 sg13g2_fill_8 FILLER_0_85_842 ();
 sg13g2_fill_1 FILLER_0_85_850 ();
 sg13g2_fill_8 FILLER_0_85_857 ();
 sg13g2_fill_4 FILLER_0_85_865 ();
 sg13g2_fill_2 FILLER_0_85_869 ();
 sg13g2_fill_1 FILLER_0_85_871 ();
 sg13g2_fill_8 FILLER_0_85_876 ();
 sg13g2_fill_8 FILLER_0_85_884 ();
 sg13g2_fill_8 FILLER_0_85_892 ();
 sg13g2_fill_8 FILLER_0_85_900 ();
 sg13g2_fill_4 FILLER_0_85_908 ();
 sg13g2_fill_4 FILLER_0_85_916 ();
 sg13g2_fill_2 FILLER_0_85_920 ();
 sg13g2_fill_1 FILLER_0_85_922 ();
 sg13g2_fill_4 FILLER_0_85_927 ();
 sg13g2_fill_1 FILLER_0_85_931 ();
 sg13g2_fill_2 FILLER_0_85_937 ();
 sg13g2_fill_2 FILLER_0_85_945 ();
 sg13g2_fill_2 FILLER_0_85_952 ();
 sg13g2_fill_8 FILLER_0_85_959 ();
 sg13g2_fill_1 FILLER_0_85_967 ();
 sg13g2_fill_8 FILLER_0_85_972 ();
 sg13g2_fill_1 FILLER_0_85_980 ();
 sg13g2_fill_2 FILLER_0_85_986 ();
 sg13g2_fill_2 FILLER_0_85_993 ();
 sg13g2_fill_8 FILLER_0_85_1000 ();
 sg13g2_fill_1 FILLER_0_85_1008 ();
 sg13g2_fill_2 FILLER_0_85_1013 ();
 sg13g2_fill_4 FILLER_0_85_1019 ();
 sg13g2_fill_2 FILLER_0_85_1023 ();
 sg13g2_fill_4 FILLER_0_85_1030 ();
 sg13g2_fill_2 FILLER_0_85_1034 ();
 sg13g2_fill_4 FILLER_0_85_1040 ();
 sg13g2_fill_2 FILLER_0_85_1044 ();
 sg13g2_fill_1 FILLER_0_85_1046 ();
 sg13g2_fill_8 FILLER_0_85_1053 ();
 sg13g2_fill_8 FILLER_0_85_1061 ();
 sg13g2_fill_2 FILLER_0_85_1069 ();
 sg13g2_fill_8 FILLER_0_85_1076 ();
 sg13g2_fill_8 FILLER_0_85_1084 ();
 sg13g2_fill_8 FILLER_0_85_1092 ();
 sg13g2_fill_8 FILLER_0_85_1100 ();
 sg13g2_fill_8 FILLER_0_85_1108 ();
 sg13g2_fill_8 FILLER_0_85_1116 ();
 sg13g2_fill_8 FILLER_0_85_1124 ();
 sg13g2_fill_4 FILLER_0_85_1132 ();
 sg13g2_fill_2 FILLER_0_85_1140 ();
 sg13g2_fill_2 FILLER_0_85_1147 ();
 sg13g2_fill_2 FILLER_0_85_1154 ();
 sg13g2_fill_2 FILLER_0_85_1161 ();
 sg13g2_fill_4 FILLER_0_85_1168 ();
 sg13g2_fill_2 FILLER_0_85_1172 ();
 sg13g2_fill_8 FILLER_0_85_1178 ();
 sg13g2_fill_4 FILLER_0_85_1191 ();
 sg13g2_fill_1 FILLER_0_85_1195 ();
 sg13g2_fill_8 FILLER_0_85_1201 ();
 sg13g2_fill_8 FILLER_0_85_1209 ();
 sg13g2_fill_8 FILLER_0_85_1217 ();
 sg13g2_fill_4 FILLER_0_85_1225 ();
 sg13g2_fill_2 FILLER_0_85_1229 ();
 sg13g2_fill_1 FILLER_0_85_1231 ();
 sg13g2_fill_8 FILLER_0_85_1237 ();
 sg13g2_fill_1 FILLER_0_85_1245 ();
 sg13g2_fill_4 FILLER_0_85_1250 ();
 sg13g2_fill_2 FILLER_0_85_1254 ();
 sg13g2_fill_1 FILLER_0_85_1256 ();
 sg13g2_fill_2 FILLER_0_85_1262 ();
 sg13g2_fill_1 FILLER_0_85_1264 ();
 sg13g2_fill_8 FILLER_0_85_1270 ();
 sg13g2_fill_2 FILLER_0_85_1283 ();
 sg13g2_fill_2 FILLER_0_85_1290 ();
 sg13g2_fill_1 FILLER_0_85_1296 ();
 sg13g2_fill_8 FILLER_0_86_0 ();
 sg13g2_fill_8 FILLER_0_86_8 ();
 sg13g2_fill_8 FILLER_0_86_16 ();
 sg13g2_fill_8 FILLER_0_86_24 ();
 sg13g2_fill_8 FILLER_0_86_32 ();
 sg13g2_fill_8 FILLER_0_86_40 ();
 sg13g2_fill_8 FILLER_0_86_48 ();
 sg13g2_fill_8 FILLER_0_86_56 ();
 sg13g2_fill_8 FILLER_0_86_64 ();
 sg13g2_fill_8 FILLER_0_86_72 ();
 sg13g2_fill_8 FILLER_0_86_80 ();
 sg13g2_fill_8 FILLER_0_86_88 ();
 sg13g2_fill_8 FILLER_0_86_96 ();
 sg13g2_fill_8 FILLER_0_86_104 ();
 sg13g2_fill_8 FILLER_0_86_112 ();
 sg13g2_fill_8 FILLER_0_86_120 ();
 sg13g2_fill_8 FILLER_0_86_128 ();
 sg13g2_fill_8 FILLER_0_86_136 ();
 sg13g2_fill_8 FILLER_0_86_144 ();
 sg13g2_fill_8 FILLER_0_86_152 ();
 sg13g2_fill_8 FILLER_0_86_160 ();
 sg13g2_fill_8 FILLER_0_86_168 ();
 sg13g2_fill_8 FILLER_0_86_176 ();
 sg13g2_fill_8 FILLER_0_86_184 ();
 sg13g2_fill_8 FILLER_0_86_192 ();
 sg13g2_fill_2 FILLER_0_86_200 ();
 sg13g2_fill_1 FILLER_0_86_202 ();
 sg13g2_fill_4 FILLER_0_86_229 ();
 sg13g2_fill_4 FILLER_0_86_254 ();
 sg13g2_fill_2 FILLER_0_86_264 ();
 sg13g2_fill_2 FILLER_0_86_292 ();
 sg13g2_fill_1 FILLER_0_86_294 ();
 sg13g2_fill_2 FILLER_0_86_299 ();
 sg13g2_fill_4 FILLER_0_86_327 ();
 sg13g2_fill_4 FILLER_0_86_336 ();
 sg13g2_fill_4 FILLER_0_86_345 ();
 sg13g2_fill_1 FILLER_0_86_349 ();
 sg13g2_fill_8 FILLER_0_86_356 ();
 sg13g2_fill_1 FILLER_0_86_364 ();
 sg13g2_fill_8 FILLER_0_86_370 ();
 sg13g2_fill_8 FILLER_0_86_378 ();
 sg13g2_fill_8 FILLER_0_86_386 ();
 sg13g2_fill_2 FILLER_0_86_394 ();
 sg13g2_fill_8 FILLER_0_86_401 ();
 sg13g2_fill_4 FILLER_0_86_413 ();
 sg13g2_fill_1 FILLER_0_86_417 ();
 sg13g2_fill_8 FILLER_0_86_423 ();
 sg13g2_fill_8 FILLER_0_86_431 ();
 sg13g2_fill_4 FILLER_0_86_439 ();
 sg13g2_fill_2 FILLER_0_86_443 ();
 sg13g2_fill_1 FILLER_0_86_445 ();
 sg13g2_fill_2 FILLER_0_86_472 ();
 sg13g2_fill_8 FILLER_0_86_479 ();
 sg13g2_fill_8 FILLER_0_86_492 ();
 sg13g2_fill_2 FILLER_0_86_505 ();
 sg13g2_fill_8 FILLER_0_86_511 ();
 sg13g2_fill_2 FILLER_0_86_519 ();
 sg13g2_fill_4 FILLER_0_86_526 ();
 sg13g2_fill_8 FILLER_0_86_534 ();
 sg13g2_fill_1 FILLER_0_86_542 ();
 sg13g2_fill_8 FILLER_0_86_548 ();
 sg13g2_fill_2 FILLER_0_86_556 ();
 sg13g2_fill_1 FILLER_0_86_558 ();
 sg13g2_fill_2 FILLER_0_86_585 ();
 sg13g2_fill_8 FILLER_0_86_592 ();
 sg13g2_fill_4 FILLER_0_86_600 ();
 sg13g2_fill_1 FILLER_0_86_604 ();
 sg13g2_fill_2 FILLER_0_86_610 ();
 sg13g2_fill_8 FILLER_0_86_616 ();
 sg13g2_fill_4 FILLER_0_86_624 ();
 sg13g2_fill_2 FILLER_0_86_628 ();
 sg13g2_fill_2 FILLER_0_86_640 ();
 sg13g2_fill_2 FILLER_0_86_647 ();
 sg13g2_fill_8 FILLER_0_86_653 ();
 sg13g2_fill_8 FILLER_0_86_661 ();
 sg13g2_fill_8 FILLER_0_86_669 ();
 sg13g2_fill_8 FILLER_0_86_677 ();
 sg13g2_fill_8 FILLER_0_86_685 ();
 sg13g2_fill_8 FILLER_0_86_693 ();
 sg13g2_fill_8 FILLER_0_86_701 ();
 sg13g2_fill_8 FILLER_0_86_709 ();
 sg13g2_fill_8 FILLER_0_86_717 ();
 sg13g2_fill_8 FILLER_0_86_725 ();
 sg13g2_fill_8 FILLER_0_86_733 ();
 sg13g2_fill_8 FILLER_0_86_741 ();
 sg13g2_fill_2 FILLER_0_86_749 ();
 sg13g2_fill_8 FILLER_0_86_757 ();
 sg13g2_fill_1 FILLER_0_86_765 ();
 sg13g2_fill_8 FILLER_0_86_770 ();
 sg13g2_fill_8 FILLER_0_86_778 ();
 sg13g2_fill_2 FILLER_0_86_786 ();
 sg13g2_fill_8 FILLER_0_86_794 ();
 sg13g2_fill_8 FILLER_0_86_802 ();
 sg13g2_fill_8 FILLER_0_86_810 ();
 sg13g2_fill_8 FILLER_0_86_818 ();
 sg13g2_fill_2 FILLER_0_86_826 ();
 sg13g2_fill_1 FILLER_0_86_828 ();
 sg13g2_fill_2 FILLER_0_86_833 ();
 sg13g2_fill_8 FILLER_0_86_840 ();
 sg13g2_fill_4 FILLER_0_86_848 ();
 sg13g2_fill_1 FILLER_0_86_852 ();
 sg13g2_fill_2 FILLER_0_86_859 ();
 sg13g2_fill_2 FILLER_0_86_867 ();
 sg13g2_fill_1 FILLER_0_86_869 ();
 sg13g2_fill_8 FILLER_0_86_878 ();
 sg13g2_fill_8 FILLER_0_86_886 ();
 sg13g2_fill_8 FILLER_0_86_894 ();
 sg13g2_fill_4 FILLER_0_86_902 ();
 sg13g2_fill_4 FILLER_0_86_910 ();
 sg13g2_fill_1 FILLER_0_86_914 ();
 sg13g2_fill_8 FILLER_0_86_921 ();
 sg13g2_fill_8 FILLER_0_86_929 ();
 sg13g2_fill_8 FILLER_0_86_942 ();
 sg13g2_fill_2 FILLER_0_86_950 ();
 sg13g2_fill_8 FILLER_0_86_957 ();
 sg13g2_fill_1 FILLER_0_86_965 ();
 sg13g2_fill_2 FILLER_0_86_970 ();
 sg13g2_fill_2 FILLER_0_86_978 ();
 sg13g2_fill_1 FILLER_0_86_980 ();
 sg13g2_fill_2 FILLER_0_86_991 ();
 sg13g2_fill_8 FILLER_0_86_997 ();
 sg13g2_fill_1 FILLER_0_86_1005 ();
 sg13g2_fill_2 FILLER_0_86_1011 ();
 sg13g2_fill_2 FILLER_0_86_1017 ();
 sg13g2_fill_1 FILLER_0_86_1019 ();
 sg13g2_fill_4 FILLER_0_86_1025 ();
 sg13g2_fill_2 FILLER_0_86_1029 ();
 sg13g2_fill_8 FILLER_0_86_1036 ();
 sg13g2_fill_4 FILLER_0_86_1044 ();
 sg13g2_fill_1 FILLER_0_86_1048 ();
 sg13g2_fill_8 FILLER_0_86_1054 ();
 sg13g2_fill_8 FILLER_0_86_1062 ();
 sg13g2_fill_8 FILLER_0_86_1070 ();
 sg13g2_fill_2 FILLER_0_86_1078 ();
 sg13g2_fill_1 FILLER_0_86_1080 ();
 sg13g2_fill_8 FILLER_0_86_1085 ();
 sg13g2_fill_8 FILLER_0_86_1093 ();
 sg13g2_fill_4 FILLER_0_86_1101 ();
 sg13g2_fill_2 FILLER_0_86_1113 ();
 sg13g2_fill_1 FILLER_0_86_1115 ();
 sg13g2_fill_2 FILLER_0_86_1121 ();
 sg13g2_fill_2 FILLER_0_86_1129 ();
 sg13g2_fill_1 FILLER_0_86_1131 ();
 sg13g2_fill_8 FILLER_0_86_1136 ();
 sg13g2_fill_8 FILLER_0_86_1144 ();
 sg13g2_fill_4 FILLER_0_86_1152 ();
 sg13g2_fill_2 FILLER_0_86_1161 ();
 sg13g2_fill_1 FILLER_0_86_1163 ();
 sg13g2_fill_8 FILLER_0_86_1169 ();
 sg13g2_fill_8 FILLER_0_86_1181 ();
 sg13g2_fill_8 FILLER_0_86_1189 ();
 sg13g2_fill_4 FILLER_0_86_1197 ();
 sg13g2_fill_4 FILLER_0_86_1204 ();
 sg13g2_fill_4 FILLER_0_86_1214 ();
 sg13g2_fill_2 FILLER_0_86_1218 ();
 sg13g2_fill_8 FILLER_0_86_1224 ();
 sg13g2_fill_8 FILLER_0_86_1232 ();
 sg13g2_fill_8 FILLER_0_86_1240 ();
 sg13g2_fill_1 FILLER_0_86_1248 ();
 sg13g2_fill_2 FILLER_0_86_1254 ();
 sg13g2_fill_8 FILLER_0_86_1260 ();
 sg13g2_fill_4 FILLER_0_86_1268 ();
 sg13g2_fill_2 FILLER_0_86_1276 ();
 sg13g2_fill_4 FILLER_0_86_1283 ();
 sg13g2_fill_1 FILLER_0_86_1287 ();
 sg13g2_fill_4 FILLER_0_86_1292 ();
 sg13g2_fill_1 FILLER_0_86_1296 ();
 sg13g2_fill_8 FILLER_0_87_0 ();
 sg13g2_fill_8 FILLER_0_87_8 ();
 sg13g2_fill_8 FILLER_0_87_16 ();
 sg13g2_fill_8 FILLER_0_87_24 ();
 sg13g2_fill_8 FILLER_0_87_32 ();
 sg13g2_fill_8 FILLER_0_87_40 ();
 sg13g2_fill_8 FILLER_0_87_48 ();
 sg13g2_fill_8 FILLER_0_87_56 ();
 sg13g2_fill_8 FILLER_0_87_64 ();
 sg13g2_fill_8 FILLER_0_87_72 ();
 sg13g2_fill_8 FILLER_0_87_80 ();
 sg13g2_fill_8 FILLER_0_87_88 ();
 sg13g2_fill_8 FILLER_0_87_96 ();
 sg13g2_fill_8 FILLER_0_87_104 ();
 sg13g2_fill_8 FILLER_0_87_112 ();
 sg13g2_fill_8 FILLER_0_87_120 ();
 sg13g2_fill_8 FILLER_0_87_128 ();
 sg13g2_fill_8 FILLER_0_87_136 ();
 sg13g2_fill_8 FILLER_0_87_144 ();
 sg13g2_fill_8 FILLER_0_87_152 ();
 sg13g2_fill_8 FILLER_0_87_160 ();
 sg13g2_fill_8 FILLER_0_87_168 ();
 sg13g2_fill_8 FILLER_0_87_176 ();
 sg13g2_fill_8 FILLER_0_87_184 ();
 sg13g2_fill_8 FILLER_0_87_192 ();
 sg13g2_fill_8 FILLER_0_87_200 ();
 sg13g2_fill_8 FILLER_0_87_208 ();
 sg13g2_fill_4 FILLER_0_87_216 ();
 sg13g2_fill_2 FILLER_0_87_220 ();
 sg13g2_fill_1 FILLER_0_87_222 ();
 sg13g2_fill_2 FILLER_0_87_228 ();
 sg13g2_fill_4 FILLER_0_87_234 ();
 sg13g2_fill_2 FILLER_0_87_238 ();
 sg13g2_fill_8 FILLER_0_87_266 ();
 sg13g2_fill_1 FILLER_0_87_274 ();
 sg13g2_fill_2 FILLER_0_87_280 ();
 sg13g2_fill_4 FILLER_0_87_287 ();
 sg13g2_fill_1 FILLER_0_87_291 ();
 sg13g2_fill_8 FILLER_0_87_296 ();
 sg13g2_fill_4 FILLER_0_87_304 ();
 sg13g2_fill_2 FILLER_0_87_308 ();
 sg13g2_fill_1 FILLER_0_87_310 ();
 sg13g2_fill_8 FILLER_0_87_316 ();
 sg13g2_fill_2 FILLER_0_87_324 ();
 sg13g2_fill_2 FILLER_0_87_331 ();
 sg13g2_fill_4 FILLER_0_87_337 ();
 sg13g2_fill_1 FILLER_0_87_341 ();
 sg13g2_fill_8 FILLER_0_87_348 ();
 sg13g2_fill_1 FILLER_0_87_356 ();
 sg13g2_fill_2 FILLER_0_87_362 ();
 sg13g2_fill_8 FILLER_0_87_368 ();
 sg13g2_fill_8 FILLER_0_87_376 ();
 sg13g2_fill_8 FILLER_0_87_384 ();
 sg13g2_fill_8 FILLER_0_87_392 ();
 sg13g2_fill_8 FILLER_0_87_407 ();
 sg13g2_fill_1 FILLER_0_87_415 ();
 sg13g2_fill_2 FILLER_0_87_421 ();
 sg13g2_fill_2 FILLER_0_87_433 ();
 sg13g2_fill_2 FILLER_0_87_440 ();
 sg13g2_fill_8 FILLER_0_87_448 ();
 sg13g2_fill_8 FILLER_0_87_456 ();
 sg13g2_fill_2 FILLER_0_87_469 ();
 sg13g2_fill_4 FILLER_0_87_475 ();
 sg13g2_fill_2 FILLER_0_87_479 ();
 sg13g2_fill_1 FILLER_0_87_481 ();
 sg13g2_fill_2 FILLER_0_87_508 ();
 sg13g2_fill_1 FILLER_0_87_510 ();
 sg13g2_fill_2 FILLER_0_87_537 ();
 sg13g2_fill_8 FILLER_0_87_549 ();
 sg13g2_fill_4 FILLER_0_87_557 ();
 sg13g2_fill_4 FILLER_0_87_582 ();
 sg13g2_fill_1 FILLER_0_87_586 ();
 sg13g2_fill_8 FILLER_0_87_591 ();
 sg13g2_fill_8 FILLER_0_87_599 ();
 sg13g2_fill_8 FILLER_0_87_607 ();
 sg13g2_fill_4 FILLER_0_87_615 ();
 sg13g2_fill_2 FILLER_0_87_619 ();
 sg13g2_fill_1 FILLER_0_87_621 ();
 sg13g2_fill_2 FILLER_0_87_627 ();
 sg13g2_fill_8 FILLER_0_87_655 ();
 sg13g2_fill_8 FILLER_0_87_663 ();
 sg13g2_fill_8 FILLER_0_87_671 ();
 sg13g2_fill_8 FILLER_0_87_679 ();
 sg13g2_fill_8 FILLER_0_87_687 ();
 sg13g2_fill_1 FILLER_0_87_695 ();
 sg13g2_fill_4 FILLER_0_87_706 ();
 sg13g2_fill_2 FILLER_0_87_710 ();
 sg13g2_fill_1 FILLER_0_87_712 ();
 sg13g2_fill_4 FILLER_0_87_717 ();
 sg13g2_fill_2 FILLER_0_87_721 ();
 sg13g2_fill_1 FILLER_0_87_723 ();
 sg13g2_fill_8 FILLER_0_87_734 ();
 sg13g2_fill_2 FILLER_0_87_742 ();
 sg13g2_fill_1 FILLER_0_87_744 ();
 sg13g2_fill_4 FILLER_0_87_749 ();
 sg13g2_fill_2 FILLER_0_87_753 ();
 sg13g2_fill_8 FILLER_0_87_765 ();
 sg13g2_fill_2 FILLER_0_87_773 ();
 sg13g2_fill_1 FILLER_0_87_775 ();
 sg13g2_fill_2 FILLER_0_87_781 ();
 sg13g2_fill_4 FILLER_0_87_789 ();
 sg13g2_fill_2 FILLER_0_87_793 ();
 sg13g2_fill_8 FILLER_0_87_805 ();
 sg13g2_fill_8 FILLER_0_87_813 ();
 sg13g2_fill_4 FILLER_0_87_821 ();
 sg13g2_fill_2 FILLER_0_87_825 ();
 sg13g2_fill_2 FILLER_0_87_834 ();
 sg13g2_fill_4 FILLER_0_87_840 ();
 sg13g2_fill_4 FILLER_0_87_850 ();
 sg13g2_fill_1 FILLER_0_87_854 ();
 sg13g2_fill_4 FILLER_0_87_859 ();
 sg13g2_fill_1 FILLER_0_87_863 ();
 sg13g2_fill_4 FILLER_0_87_868 ();
 sg13g2_fill_1 FILLER_0_87_872 ();
 sg13g2_fill_8 FILLER_0_87_880 ();
 sg13g2_fill_8 FILLER_0_87_888 ();
 sg13g2_fill_8 FILLER_0_87_896 ();
 sg13g2_fill_8 FILLER_0_87_904 ();
 sg13g2_fill_4 FILLER_0_87_912 ();
 sg13g2_fill_2 FILLER_0_87_916 ();
 sg13g2_fill_2 FILLER_0_87_924 ();
 sg13g2_fill_4 FILLER_0_87_931 ();
 sg13g2_fill_2 FILLER_0_87_935 ();
 sg13g2_fill_8 FILLER_0_87_941 ();
 sg13g2_fill_8 FILLER_0_87_949 ();
 sg13g2_fill_8 FILLER_0_87_957 ();
 sg13g2_fill_8 FILLER_0_87_965 ();
 sg13g2_fill_1 FILLER_0_87_973 ();
 sg13g2_fill_2 FILLER_0_87_979 ();
 sg13g2_fill_8 FILLER_0_87_986 ();
 sg13g2_fill_1 FILLER_0_87_994 ();
 sg13g2_fill_8 FILLER_0_87_999 ();
 sg13g2_fill_1 FILLER_0_87_1007 ();
 sg13g2_fill_4 FILLER_0_87_1012 ();
 sg13g2_fill_1 FILLER_0_87_1016 ();
 sg13g2_fill_2 FILLER_0_87_1023 ();
 sg13g2_fill_2 FILLER_0_87_1030 ();
 sg13g2_fill_2 FILLER_0_87_1038 ();
 sg13g2_fill_8 FILLER_0_87_1046 ();
 sg13g2_fill_8 FILLER_0_87_1054 ();
 sg13g2_fill_8 FILLER_0_87_1062 ();
 sg13g2_fill_8 FILLER_0_87_1070 ();
 sg13g2_fill_8 FILLER_0_87_1078 ();
 sg13g2_fill_8 FILLER_0_87_1086 ();
 sg13g2_fill_8 FILLER_0_87_1094 ();
 sg13g2_fill_8 FILLER_0_87_1102 ();
 sg13g2_fill_8 FILLER_0_87_1110 ();
 sg13g2_fill_4 FILLER_0_87_1118 ();
 sg13g2_fill_8 FILLER_0_87_1128 ();
 sg13g2_fill_8 FILLER_0_87_1136 ();
 sg13g2_fill_2 FILLER_0_87_1149 ();
 sg13g2_fill_8 FILLER_0_87_1156 ();
 sg13g2_fill_4 FILLER_0_87_1164 ();
 sg13g2_fill_2 FILLER_0_87_1168 ();
 sg13g2_fill_8 FILLER_0_87_1175 ();
 sg13g2_fill_1 FILLER_0_87_1183 ();
 sg13g2_fill_2 FILLER_0_87_1191 ();
 sg13g2_fill_4 FILLER_0_87_1198 ();
 sg13g2_fill_2 FILLER_0_87_1208 ();
 sg13g2_fill_1 FILLER_0_87_1210 ();
 sg13g2_fill_2 FILLER_0_87_1217 ();
 sg13g2_fill_1 FILLER_0_87_1219 ();
 sg13g2_fill_2 FILLER_0_87_1227 ();
 sg13g2_fill_2 FILLER_0_87_1236 ();
 sg13g2_fill_2 FILLER_0_87_1244 ();
 sg13g2_fill_4 FILLER_0_87_1250 ();
 sg13g2_fill_2 FILLER_0_87_1254 ();
 sg13g2_fill_1 FILLER_0_87_1256 ();
 sg13g2_fill_8 FILLER_0_87_1262 ();
 sg13g2_fill_1 FILLER_0_87_1270 ();
 sg13g2_fill_2 FILLER_0_87_1276 ();
 sg13g2_fill_4 FILLER_0_87_1286 ();
 sg13g2_fill_2 FILLER_0_87_1294 ();
 sg13g2_fill_1 FILLER_0_87_1296 ();
 sg13g2_fill_8 FILLER_0_88_0 ();
 sg13g2_fill_8 FILLER_0_88_8 ();
 sg13g2_fill_8 FILLER_0_88_16 ();
 sg13g2_fill_8 FILLER_0_88_24 ();
 sg13g2_fill_8 FILLER_0_88_32 ();
 sg13g2_fill_8 FILLER_0_88_40 ();
 sg13g2_fill_8 FILLER_0_88_48 ();
 sg13g2_fill_8 FILLER_0_88_56 ();
 sg13g2_fill_8 FILLER_0_88_64 ();
 sg13g2_fill_8 FILLER_0_88_72 ();
 sg13g2_fill_8 FILLER_0_88_80 ();
 sg13g2_fill_8 FILLER_0_88_88 ();
 sg13g2_fill_8 FILLER_0_88_96 ();
 sg13g2_fill_8 FILLER_0_88_104 ();
 sg13g2_fill_8 FILLER_0_88_112 ();
 sg13g2_fill_8 FILLER_0_88_120 ();
 sg13g2_fill_8 FILLER_0_88_128 ();
 sg13g2_fill_8 FILLER_0_88_136 ();
 sg13g2_fill_8 FILLER_0_88_144 ();
 sg13g2_fill_8 FILLER_0_88_152 ();
 sg13g2_fill_8 FILLER_0_88_160 ();
 sg13g2_fill_8 FILLER_0_88_168 ();
 sg13g2_fill_8 FILLER_0_88_176 ();
 sg13g2_fill_8 FILLER_0_88_184 ();
 sg13g2_fill_8 FILLER_0_88_192 ();
 sg13g2_fill_8 FILLER_0_88_200 ();
 sg13g2_fill_8 FILLER_0_88_208 ();
 sg13g2_fill_2 FILLER_0_88_242 ();
 sg13g2_fill_2 FILLER_0_88_249 ();
 sg13g2_fill_2 FILLER_0_88_255 ();
 sg13g2_fill_8 FILLER_0_88_262 ();
 sg13g2_fill_8 FILLER_0_88_270 ();
 sg13g2_fill_8 FILLER_0_88_278 ();
 sg13g2_fill_8 FILLER_0_88_286 ();
 sg13g2_fill_8 FILLER_0_88_294 ();
 sg13g2_fill_8 FILLER_0_88_302 ();
 sg13g2_fill_8 FILLER_0_88_310 ();
 sg13g2_fill_4 FILLER_0_88_318 ();
 sg13g2_fill_1 FILLER_0_88_322 ();
 sg13g2_fill_4 FILLER_0_88_349 ();
 sg13g2_fill_2 FILLER_0_88_353 ();
 sg13g2_fill_8 FILLER_0_88_381 ();
 sg13g2_fill_8 FILLER_0_88_389 ();
 sg13g2_fill_2 FILLER_0_88_397 ();
 sg13g2_fill_2 FILLER_0_88_405 ();
 sg13g2_fill_1 FILLER_0_88_407 ();
 sg13g2_fill_2 FILLER_0_88_413 ();
 sg13g2_fill_4 FILLER_0_88_419 ();
 sg13g2_fill_2 FILLER_0_88_427 ();
 sg13g2_fill_1 FILLER_0_88_429 ();
 sg13g2_fill_8 FILLER_0_88_456 ();
 sg13g2_fill_8 FILLER_0_88_464 ();
 sg13g2_fill_8 FILLER_0_88_472 ();
 sg13g2_fill_4 FILLER_0_88_480 ();
 sg13g2_fill_1 FILLER_0_88_484 ();
 sg13g2_fill_8 FILLER_0_88_489 ();
 sg13g2_fill_2 FILLER_0_88_502 ();
 sg13g2_fill_8 FILLER_0_88_510 ();
 sg13g2_fill_8 FILLER_0_88_518 ();
 sg13g2_fill_8 FILLER_0_88_526 ();
 sg13g2_fill_8 FILLER_0_88_534 ();
 sg13g2_fill_8 FILLER_0_88_542 ();
 sg13g2_fill_8 FILLER_0_88_550 ();
 sg13g2_fill_4 FILLER_0_88_558 ();
 sg13g2_fill_2 FILLER_0_88_562 ();
 sg13g2_fill_1 FILLER_0_88_564 ();
 sg13g2_fill_8 FILLER_0_88_575 ();
 sg13g2_fill_8 FILLER_0_88_583 ();
 sg13g2_fill_8 FILLER_0_88_591 ();
 sg13g2_fill_4 FILLER_0_88_599 ();
 sg13g2_fill_2 FILLER_0_88_603 ();
 sg13g2_fill_1 FILLER_0_88_605 ();
 sg13g2_fill_4 FILLER_0_88_632 ();
 sg13g2_fill_2 FILLER_0_88_636 ();
 sg13g2_fill_2 FILLER_0_88_643 ();
 sg13g2_fill_2 FILLER_0_88_650 ();
 sg13g2_fill_4 FILLER_0_88_657 ();
 sg13g2_fill_2 FILLER_0_88_671 ();
 sg13g2_fill_1 FILLER_0_88_673 ();
 sg13g2_fill_2 FILLER_0_88_700 ();
 sg13g2_fill_1 FILLER_0_88_702 ();
 sg13g2_fill_2 FILLER_0_88_729 ();
 sg13g2_fill_2 FILLER_0_88_757 ();
 sg13g2_fill_2 FILLER_0_88_785 ();
 sg13g2_fill_4 FILLER_0_88_813 ();
 sg13g2_fill_8 FILLER_0_88_821 ();
 sg13g2_fill_2 FILLER_0_88_834 ();
 sg13g2_fill_8 FILLER_0_88_841 ();
 sg13g2_fill_2 FILLER_0_88_853 ();
 sg13g2_fill_2 FILLER_0_88_864 ();
 sg13g2_fill_2 FILLER_0_88_872 ();
 sg13g2_fill_2 FILLER_0_88_878 ();
 sg13g2_fill_2 FILLER_0_88_885 ();
 sg13g2_fill_1 FILLER_0_88_887 ();
 sg13g2_fill_8 FILLER_0_88_894 ();
 sg13g2_fill_8 FILLER_0_88_905 ();
 sg13g2_fill_2 FILLER_0_88_913 ();
 sg13g2_fill_1 FILLER_0_88_915 ();
 sg13g2_fill_8 FILLER_0_88_921 ();
 sg13g2_fill_8 FILLER_0_88_929 ();
 sg13g2_fill_2 FILLER_0_88_937 ();
 sg13g2_fill_2 FILLER_0_88_944 ();
 sg13g2_fill_2 FILLER_0_88_951 ();
 sg13g2_fill_2 FILLER_0_88_957 ();
 sg13g2_fill_1 FILLER_0_88_959 ();
 sg13g2_fill_8 FILLER_0_88_964 ();
 sg13g2_fill_8 FILLER_0_88_972 ();
 sg13g2_fill_4 FILLER_0_88_980 ();
 sg13g2_fill_2 FILLER_0_88_988 ();
 sg13g2_fill_2 FILLER_0_88_994 ();
 sg13g2_fill_1 FILLER_0_88_996 ();
 sg13g2_fill_8 FILLER_0_88_1002 ();
 sg13g2_fill_2 FILLER_0_88_1010 ();
 sg13g2_fill_2 FILLER_0_88_1017 ();
 sg13g2_fill_2 FILLER_0_88_1023 ();
 sg13g2_fill_2 FILLER_0_88_1030 ();
 sg13g2_fill_2 FILLER_0_88_1037 ();
 sg13g2_fill_8 FILLER_0_88_1043 ();
 sg13g2_fill_8 FILLER_0_88_1051 ();
 sg13g2_fill_8 FILLER_0_88_1059 ();
 sg13g2_fill_4 FILLER_0_88_1072 ();
 sg13g2_fill_1 FILLER_0_88_1076 ();
 sg13g2_fill_2 FILLER_0_88_1083 ();
 sg13g2_fill_8 FILLER_0_88_1089 ();
 sg13g2_fill_1 FILLER_0_88_1097 ();
 sg13g2_fill_2 FILLER_0_88_1105 ();
 sg13g2_fill_2 FILLER_0_88_1112 ();
 sg13g2_fill_2 FILLER_0_88_1119 ();
 sg13g2_fill_2 FILLER_0_88_1126 ();
 sg13g2_fill_2 FILLER_0_88_1132 ();
 sg13g2_fill_1 FILLER_0_88_1134 ();
 sg13g2_fill_2 FILLER_0_88_1147 ();
 sg13g2_fill_2 FILLER_0_88_1157 ();
 sg13g2_fill_2 FILLER_0_88_1164 ();
 sg13g2_fill_1 FILLER_0_88_1166 ();
 sg13g2_fill_2 FILLER_0_88_1170 ();
 sg13g2_fill_4 FILLER_0_88_1178 ();
 sg13g2_fill_8 FILLER_0_88_1186 ();
 sg13g2_fill_2 FILLER_0_88_1194 ();
 sg13g2_fill_4 FILLER_0_88_1203 ();
 sg13g2_fill_2 FILLER_0_88_1215 ();
 sg13g2_fill_1 FILLER_0_88_1217 ();
 sg13g2_fill_2 FILLER_0_88_1225 ();
 sg13g2_fill_8 FILLER_0_88_1231 ();
 sg13g2_fill_4 FILLER_0_88_1239 ();
 sg13g2_fill_2 FILLER_0_88_1247 ();
 sg13g2_fill_2 FILLER_0_88_1253 ();
 sg13g2_fill_8 FILLER_0_88_1263 ();
 sg13g2_fill_2 FILLER_0_88_1271 ();
 sg13g2_fill_1 FILLER_0_88_1273 ();
 sg13g2_fill_2 FILLER_0_88_1278 ();
 sg13g2_fill_2 FILLER_0_88_1283 ();
 sg13g2_fill_8 FILLER_0_88_1289 ();
 sg13g2_fill_8 FILLER_0_89_0 ();
 sg13g2_fill_8 FILLER_0_89_8 ();
 sg13g2_fill_8 FILLER_0_89_16 ();
 sg13g2_fill_8 FILLER_0_89_24 ();
 sg13g2_fill_8 FILLER_0_89_32 ();
 sg13g2_fill_8 FILLER_0_89_40 ();
 sg13g2_fill_8 FILLER_0_89_48 ();
 sg13g2_fill_8 FILLER_0_89_56 ();
 sg13g2_fill_8 FILLER_0_89_64 ();
 sg13g2_fill_8 FILLER_0_89_72 ();
 sg13g2_fill_8 FILLER_0_89_80 ();
 sg13g2_fill_8 FILLER_0_89_88 ();
 sg13g2_fill_8 FILLER_0_89_96 ();
 sg13g2_fill_8 FILLER_0_89_104 ();
 sg13g2_fill_8 FILLER_0_89_112 ();
 sg13g2_fill_8 FILLER_0_89_120 ();
 sg13g2_fill_8 FILLER_0_89_128 ();
 sg13g2_fill_8 FILLER_0_89_136 ();
 sg13g2_fill_8 FILLER_0_89_144 ();
 sg13g2_fill_8 FILLER_0_89_152 ();
 sg13g2_fill_8 FILLER_0_89_160 ();
 sg13g2_fill_8 FILLER_0_89_168 ();
 sg13g2_fill_8 FILLER_0_89_176 ();
 sg13g2_fill_8 FILLER_0_89_184 ();
 sg13g2_fill_8 FILLER_0_89_192 ();
 sg13g2_fill_8 FILLER_0_89_200 ();
 sg13g2_fill_2 FILLER_0_89_208 ();
 sg13g2_fill_1 FILLER_0_89_210 ();
 sg13g2_fill_8 FILLER_0_89_216 ();
 sg13g2_fill_8 FILLER_0_89_228 ();
 sg13g2_fill_8 FILLER_0_89_236 ();
 sg13g2_fill_8 FILLER_0_89_244 ();
 sg13g2_fill_8 FILLER_0_89_252 ();
 sg13g2_fill_1 FILLER_0_89_260 ();
 sg13g2_fill_8 FILLER_0_89_266 ();
 sg13g2_fill_8 FILLER_0_89_274 ();
 sg13g2_fill_8 FILLER_0_89_282 ();
 sg13g2_fill_8 FILLER_0_89_290 ();
 sg13g2_fill_8 FILLER_0_89_298 ();
 sg13g2_fill_8 FILLER_0_89_306 ();
 sg13g2_fill_8 FILLER_0_89_314 ();
 sg13g2_fill_8 FILLER_0_89_322 ();
 sg13g2_fill_8 FILLER_0_89_330 ();
 sg13g2_fill_8 FILLER_0_89_338 ();
 sg13g2_fill_8 FILLER_0_89_346 ();
 sg13g2_fill_4 FILLER_0_89_354 ();
 sg13g2_fill_2 FILLER_0_89_358 ();
 sg13g2_fill_4 FILLER_0_89_381 ();
 sg13g2_fill_2 FILLER_0_89_385 ();
 sg13g2_fill_1 FILLER_0_89_387 ();
 sg13g2_fill_4 FILLER_0_89_414 ();
 sg13g2_fill_1 FILLER_0_89_418 ();
 sg13g2_fill_4 FILLER_0_89_424 ();
 sg13g2_fill_4 FILLER_0_89_433 ();
 sg13g2_fill_8 FILLER_0_89_442 ();
 sg13g2_fill_8 FILLER_0_89_450 ();
 sg13g2_fill_8 FILLER_0_89_458 ();
 sg13g2_fill_8 FILLER_0_89_466 ();
 sg13g2_fill_2 FILLER_0_89_474 ();
 sg13g2_fill_1 FILLER_0_89_476 ();
 sg13g2_fill_2 FILLER_0_89_482 ();
 sg13g2_fill_2 FILLER_0_89_489 ();
 sg13g2_fill_8 FILLER_0_89_517 ();
 sg13g2_fill_8 FILLER_0_89_525 ();
 sg13g2_fill_2 FILLER_0_89_533 ();
 sg13g2_fill_1 FILLER_0_89_535 ();
 sg13g2_fill_2 FILLER_0_89_541 ();
 sg13g2_fill_2 FILLER_0_89_569 ();
 sg13g2_fill_8 FILLER_0_89_575 ();
 sg13g2_fill_4 FILLER_0_89_583 ();
 sg13g2_fill_2 FILLER_0_89_587 ();
 sg13g2_fill_4 FILLER_0_89_593 ();
 sg13g2_fill_8 FILLER_0_89_602 ();
 sg13g2_fill_8 FILLER_0_89_610 ();
 sg13g2_fill_1 FILLER_0_89_618 ();
 sg13g2_fill_8 FILLER_0_89_625 ();
 sg13g2_fill_1 FILLER_0_89_633 ();
 sg13g2_fill_8 FILLER_0_89_638 ();
 sg13g2_fill_2 FILLER_0_89_646 ();
 sg13g2_fill_2 FILLER_0_89_658 ();
 sg13g2_fill_2 FILLER_0_89_686 ();
 sg13g2_fill_2 FILLER_0_89_709 ();
 sg13g2_fill_2 FILLER_0_89_716 ();
 sg13g2_fill_1 FILLER_0_89_718 ();
 sg13g2_fill_8 FILLER_0_89_724 ();
 sg13g2_fill_8 FILLER_0_89_732 ();
 sg13g2_fill_8 FILLER_0_89_740 ();
 sg13g2_fill_8 FILLER_0_89_748 ();
 sg13g2_fill_1 FILLER_0_89_756 ();
 sg13g2_fill_8 FILLER_0_89_762 ();
 sg13g2_fill_8 FILLER_0_89_770 ();
 sg13g2_fill_1 FILLER_0_89_778 ();
 sg13g2_fill_8 FILLER_0_89_784 ();
 sg13g2_fill_8 FILLER_0_89_792 ();
 sg13g2_fill_8 FILLER_0_89_800 ();
 sg13g2_fill_8 FILLER_0_89_808 ();
 sg13g2_fill_8 FILLER_0_89_816 ();
 sg13g2_fill_4 FILLER_0_89_824 ();
 sg13g2_fill_2 FILLER_0_89_834 ();
 sg13g2_fill_2 FILLER_0_89_841 ();
 sg13g2_fill_1 FILLER_0_89_843 ();
 sg13g2_fill_2 FILLER_0_89_856 ();
 sg13g2_fill_2 FILLER_0_89_863 ();
 sg13g2_fill_2 FILLER_0_89_874 ();
 sg13g2_fill_2 FILLER_0_89_882 ();
 sg13g2_fill_8 FILLER_0_89_893 ();
 sg13g2_fill_2 FILLER_0_89_901 ();
 sg13g2_fill_1 FILLER_0_89_903 ();
 sg13g2_fill_8 FILLER_0_89_908 ();
 sg13g2_fill_4 FILLER_0_89_916 ();
 sg13g2_fill_1 FILLER_0_89_920 ();
 sg13g2_fill_4 FILLER_0_89_925 ();
 sg13g2_fill_2 FILLER_0_89_929 ();
 sg13g2_fill_2 FILLER_0_89_936 ();
 sg13g2_fill_2 FILLER_0_89_942 ();
 sg13g2_fill_4 FILLER_0_89_950 ();
 sg13g2_fill_2 FILLER_0_89_954 ();
 sg13g2_fill_1 FILLER_0_89_956 ();
 sg13g2_fill_2 FILLER_0_89_961 ();
 sg13g2_fill_4 FILLER_0_89_968 ();
 sg13g2_fill_1 FILLER_0_89_972 ();
 sg13g2_fill_2 FILLER_0_89_979 ();
 sg13g2_fill_4 FILLER_0_89_986 ();
 sg13g2_fill_2 FILLER_0_89_990 ();
 sg13g2_fill_2 FILLER_0_89_998 ();
 sg13g2_fill_1 FILLER_0_89_1000 ();
 sg13g2_fill_2 FILLER_0_89_1005 ();
 sg13g2_fill_1 FILLER_0_89_1007 ();
 sg13g2_fill_2 FILLER_0_89_1013 ();
 sg13g2_fill_2 FILLER_0_89_1019 ();
 sg13g2_fill_8 FILLER_0_89_1026 ();
 sg13g2_fill_8 FILLER_0_89_1039 ();
 sg13g2_fill_8 FILLER_0_89_1047 ();
 sg13g2_fill_4 FILLER_0_89_1055 ();
 sg13g2_fill_1 FILLER_0_89_1059 ();
 sg13g2_fill_2 FILLER_0_89_1064 ();
 sg13g2_fill_2 FILLER_0_89_1072 ();
 sg13g2_fill_2 FILLER_0_89_1079 ();
 sg13g2_fill_2 FILLER_0_89_1086 ();
 sg13g2_fill_2 FILLER_0_89_1093 ();
 sg13g2_fill_2 FILLER_0_89_1102 ();
 sg13g2_fill_2 FILLER_0_89_1110 ();
 sg13g2_fill_2 FILLER_0_89_1117 ();
 sg13g2_fill_2 FILLER_0_89_1123 ();
 sg13g2_fill_2 FILLER_0_89_1130 ();
 sg13g2_fill_2 FILLER_0_89_1137 ();
 sg13g2_fill_4 FILLER_0_89_1145 ();
 sg13g2_fill_2 FILLER_0_89_1153 ();
 sg13g2_fill_4 FILLER_0_89_1160 ();
 sg13g2_fill_1 FILLER_0_89_1164 ();
 sg13g2_fill_4 FILLER_0_89_1171 ();
 sg13g2_fill_1 FILLER_0_89_1175 ();
 sg13g2_fill_2 FILLER_0_89_1181 ();
 sg13g2_fill_4 FILLER_0_89_1188 ();
 sg13g2_fill_1 FILLER_0_89_1192 ();
 sg13g2_fill_4 FILLER_0_89_1198 ();
 sg13g2_fill_2 FILLER_0_89_1207 ();
 sg13g2_fill_2 FILLER_0_89_1214 ();
 sg13g2_fill_1 FILLER_0_89_1216 ();
 sg13g2_fill_2 FILLER_0_89_1224 ();
 sg13g2_fill_8 FILLER_0_89_1230 ();
 sg13g2_fill_8 FILLER_0_89_1238 ();
 sg13g2_fill_2 FILLER_0_89_1246 ();
 sg13g2_fill_1 FILLER_0_89_1248 ();
 sg13g2_fill_2 FILLER_0_89_1259 ();
 sg13g2_fill_2 FILLER_0_89_1266 ();
 sg13g2_fill_4 FILLER_0_89_1276 ();
 sg13g2_fill_2 FILLER_0_89_1280 ();
 sg13g2_fill_1 FILLER_0_89_1282 ();
 sg13g2_fill_8 FILLER_0_89_1288 ();
 sg13g2_fill_1 FILLER_0_89_1296 ();
 sg13g2_fill_8 FILLER_0_90_0 ();
 sg13g2_fill_8 FILLER_0_90_8 ();
 sg13g2_fill_8 FILLER_0_90_16 ();
 sg13g2_fill_8 FILLER_0_90_24 ();
 sg13g2_fill_8 FILLER_0_90_32 ();
 sg13g2_fill_8 FILLER_0_90_40 ();
 sg13g2_fill_8 FILLER_0_90_48 ();
 sg13g2_fill_8 FILLER_0_90_56 ();
 sg13g2_fill_8 FILLER_0_90_64 ();
 sg13g2_fill_8 FILLER_0_90_72 ();
 sg13g2_fill_8 FILLER_0_90_80 ();
 sg13g2_fill_8 FILLER_0_90_88 ();
 sg13g2_fill_8 FILLER_0_90_96 ();
 sg13g2_fill_8 FILLER_0_90_104 ();
 sg13g2_fill_8 FILLER_0_90_112 ();
 sg13g2_fill_8 FILLER_0_90_120 ();
 sg13g2_fill_8 FILLER_0_90_128 ();
 sg13g2_fill_8 FILLER_0_90_136 ();
 sg13g2_fill_8 FILLER_0_90_144 ();
 sg13g2_fill_8 FILLER_0_90_152 ();
 sg13g2_fill_8 FILLER_0_90_160 ();
 sg13g2_fill_8 FILLER_0_90_168 ();
 sg13g2_fill_8 FILLER_0_90_176 ();
 sg13g2_fill_8 FILLER_0_90_184 ();
 sg13g2_fill_8 FILLER_0_90_192 ();
 sg13g2_fill_8 FILLER_0_90_200 ();
 sg13g2_fill_8 FILLER_0_90_208 ();
 sg13g2_fill_8 FILLER_0_90_216 ();
 sg13g2_fill_8 FILLER_0_90_224 ();
 sg13g2_fill_8 FILLER_0_90_232 ();
 sg13g2_fill_8 FILLER_0_90_240 ();
 sg13g2_fill_8 FILLER_0_90_248 ();
 sg13g2_fill_8 FILLER_0_90_256 ();
 sg13g2_fill_1 FILLER_0_90_264 ();
 sg13g2_fill_8 FILLER_0_90_270 ();
 sg13g2_fill_8 FILLER_0_90_278 ();
 sg13g2_fill_8 FILLER_0_90_286 ();
 sg13g2_fill_8 FILLER_0_90_294 ();
 sg13g2_fill_8 FILLER_0_90_302 ();
 sg13g2_fill_8 FILLER_0_90_310 ();
 sg13g2_fill_8 FILLER_0_90_318 ();
 sg13g2_fill_8 FILLER_0_90_326 ();
 sg13g2_fill_4 FILLER_0_90_334 ();
 sg13g2_fill_4 FILLER_0_90_364 ();
 sg13g2_fill_2 FILLER_0_90_368 ();
 sg13g2_fill_8 FILLER_0_90_375 ();
 sg13g2_fill_8 FILLER_0_90_383 ();
 sg13g2_fill_1 FILLER_0_90_391 ();
 sg13g2_fill_8 FILLER_0_90_396 ();
 sg13g2_fill_8 FILLER_0_90_404 ();
 sg13g2_fill_1 FILLER_0_90_412 ();
 sg13g2_fill_4 FILLER_0_90_419 ();
 sg13g2_fill_8 FILLER_0_90_427 ();
 sg13g2_fill_8 FILLER_0_90_435 ();
 sg13g2_fill_8 FILLER_0_90_443 ();
 sg13g2_fill_1 FILLER_0_90_451 ();
 sg13g2_fill_4 FILLER_0_90_460 ();
 sg13g2_fill_2 FILLER_0_90_464 ();
 sg13g2_fill_1 FILLER_0_90_466 ();
 sg13g2_fill_2 FILLER_0_90_472 ();
 sg13g2_fill_4 FILLER_0_90_479 ();
 sg13g2_fill_1 FILLER_0_90_483 ();
 sg13g2_fill_2 FILLER_0_90_488 ();
 sg13g2_fill_2 FILLER_0_90_495 ();
 sg13g2_fill_4 FILLER_0_90_501 ();
 sg13g2_fill_2 FILLER_0_90_505 ();
 sg13g2_fill_2 FILLER_0_90_528 ();
 sg13g2_fill_2 FILLER_0_90_535 ();
 sg13g2_fill_8 FILLER_0_90_541 ();
 sg13g2_fill_8 FILLER_0_90_549 ();
 sg13g2_fill_2 FILLER_0_90_557 ();
 sg13g2_fill_2 FILLER_0_90_564 ();
 sg13g2_fill_4 FILLER_0_90_571 ();
 sg13g2_fill_2 FILLER_0_90_601 ();
 sg13g2_fill_2 FILLER_0_90_608 ();
 sg13g2_fill_2 FILLER_0_90_616 ();
 sg13g2_fill_1 FILLER_0_90_618 ();
 sg13g2_fill_2 FILLER_0_90_625 ();
 sg13g2_fill_2 FILLER_0_90_631 ();
 sg13g2_fill_2 FILLER_0_90_638 ();
 sg13g2_fill_4 FILLER_0_90_645 ();
 sg13g2_fill_2 FILLER_0_90_649 ();
 sg13g2_fill_1 FILLER_0_90_651 ();
 sg13g2_fill_8 FILLER_0_90_656 ();
 sg13g2_fill_8 FILLER_0_90_664 ();
 sg13g2_fill_8 FILLER_0_90_672 ();
 sg13g2_fill_8 FILLER_0_90_680 ();
 sg13g2_fill_8 FILLER_0_90_688 ();
 sg13g2_fill_8 FILLER_0_90_696 ();
 sg13g2_fill_8 FILLER_0_90_708 ();
 sg13g2_fill_8 FILLER_0_90_716 ();
 sg13g2_fill_8 FILLER_0_90_724 ();
 sg13g2_fill_8 FILLER_0_90_732 ();
 sg13g2_fill_4 FILLER_0_90_740 ();
 sg13g2_fill_2 FILLER_0_90_744 ();
 sg13g2_fill_1 FILLER_0_90_746 ();
 sg13g2_fill_2 FILLER_0_90_757 ();
 sg13g2_fill_2 FILLER_0_90_764 ();
 sg13g2_fill_8 FILLER_0_90_774 ();
 sg13g2_fill_8 FILLER_0_90_782 ();
 sg13g2_fill_8 FILLER_0_90_790 ();
 sg13g2_fill_4 FILLER_0_90_798 ();
 sg13g2_fill_2 FILLER_0_90_802 ();
 sg13g2_fill_1 FILLER_0_90_804 ();
 sg13g2_fill_4 FILLER_0_90_810 ();
 sg13g2_fill_1 FILLER_0_90_814 ();
 sg13g2_fill_8 FILLER_0_90_819 ();
 sg13g2_fill_2 FILLER_0_90_827 ();
 sg13g2_fill_1 FILLER_0_90_829 ();
 sg13g2_fill_4 FILLER_0_90_834 ();
 sg13g2_fill_2 FILLER_0_90_838 ();
 sg13g2_fill_1 FILLER_0_90_840 ();
 sg13g2_fill_2 FILLER_0_90_845 ();
 sg13g2_fill_8 FILLER_0_90_851 ();
 sg13g2_fill_8 FILLER_0_90_859 ();
 sg13g2_fill_8 FILLER_0_90_867 ();
 sg13g2_fill_8 FILLER_0_90_875 ();
 sg13g2_fill_8 FILLER_0_90_883 ();
 sg13g2_fill_8 FILLER_0_90_891 ();
 sg13g2_fill_8 FILLER_0_90_899 ();
 sg13g2_fill_8 FILLER_0_90_907 ();
 sg13g2_fill_2 FILLER_0_90_915 ();
 sg13g2_fill_1 FILLER_0_90_917 ();
 sg13g2_fill_4 FILLER_0_90_928 ();
 sg13g2_fill_1 FILLER_0_90_932 ();
 sg13g2_fill_8 FILLER_0_90_943 ();
 sg13g2_fill_2 FILLER_0_90_951 ();
 sg13g2_fill_1 FILLER_0_90_953 ();
 sg13g2_fill_2 FILLER_0_90_959 ();
 sg13g2_fill_8 FILLER_0_90_967 ();
 sg13g2_fill_8 FILLER_0_90_975 ();
 sg13g2_fill_4 FILLER_0_90_983 ();
 sg13g2_fill_2 FILLER_0_90_995 ();
 sg13g2_fill_4 FILLER_0_90_1000 ();
 sg13g2_fill_2 FILLER_0_90_1004 ();
 sg13g2_fill_1 FILLER_0_90_1006 ();
 sg13g2_fill_2 FILLER_0_90_1012 ();
 sg13g2_fill_2 FILLER_0_90_1020 ();
 sg13g2_fill_8 FILLER_0_90_1027 ();
 sg13g2_fill_8 FILLER_0_90_1035 ();
 sg13g2_fill_8 FILLER_0_90_1043 ();
 sg13g2_fill_4 FILLER_0_90_1051 ();
 sg13g2_fill_2 FILLER_0_90_1055 ();
 sg13g2_fill_4 FILLER_0_90_1062 ();
 sg13g2_fill_2 FILLER_0_90_1066 ();
 sg13g2_fill_1 FILLER_0_90_1068 ();
 sg13g2_fill_2 FILLER_0_90_1075 ();
 sg13g2_fill_1 FILLER_0_90_1077 ();
 sg13g2_fill_4 FILLER_0_90_1083 ();
 sg13g2_fill_2 FILLER_0_90_1087 ();
 sg13g2_fill_2 FILLER_0_90_1093 ();
 sg13g2_fill_2 FILLER_0_90_1100 ();
 sg13g2_fill_2 FILLER_0_90_1109 ();
 sg13g2_fill_2 FILLER_0_90_1115 ();
 sg13g2_fill_2 FILLER_0_90_1122 ();
 sg13g2_fill_4 FILLER_0_90_1130 ();
 sg13g2_fill_2 FILLER_0_90_1134 ();
 sg13g2_fill_8 FILLER_0_90_1140 ();
 sg13g2_fill_8 FILLER_0_90_1148 ();
 sg13g2_fill_8 FILLER_0_90_1156 ();
 sg13g2_fill_8 FILLER_0_90_1164 ();
 sg13g2_fill_8 FILLER_0_90_1177 ();
 sg13g2_fill_1 FILLER_0_90_1185 ();
 sg13g2_fill_8 FILLER_0_90_1191 ();
 sg13g2_fill_2 FILLER_0_90_1206 ();
 sg13g2_fill_2 FILLER_0_90_1213 ();
 sg13g2_fill_2 FILLER_0_90_1222 ();
 sg13g2_fill_2 FILLER_0_90_1230 ();
 sg13g2_fill_2 FILLER_0_90_1236 ();
 sg13g2_fill_1 FILLER_0_90_1238 ();
 sg13g2_fill_2 FILLER_0_90_1244 ();
 sg13g2_fill_2 FILLER_0_90_1256 ();
 sg13g2_fill_4 FILLER_0_90_1284 ();
 sg13g2_fill_2 FILLER_0_90_1288 ();
 sg13g2_fill_2 FILLER_0_90_1294 ();
 sg13g2_fill_1 FILLER_0_90_1296 ();
 sg13g2_fill_8 FILLER_0_91_0 ();
 sg13g2_fill_8 FILLER_0_91_8 ();
 sg13g2_fill_8 FILLER_0_91_16 ();
 sg13g2_fill_8 FILLER_0_91_24 ();
 sg13g2_fill_8 FILLER_0_91_32 ();
 sg13g2_fill_8 FILLER_0_91_40 ();
 sg13g2_fill_8 FILLER_0_91_48 ();
 sg13g2_fill_8 FILLER_0_91_56 ();
 sg13g2_fill_8 FILLER_0_91_64 ();
 sg13g2_fill_8 FILLER_0_91_72 ();
 sg13g2_fill_8 FILLER_0_91_80 ();
 sg13g2_fill_8 FILLER_0_91_88 ();
 sg13g2_fill_8 FILLER_0_91_96 ();
 sg13g2_fill_8 FILLER_0_91_104 ();
 sg13g2_fill_8 FILLER_0_91_112 ();
 sg13g2_fill_8 FILLER_0_91_120 ();
 sg13g2_fill_8 FILLER_0_91_128 ();
 sg13g2_fill_8 FILLER_0_91_136 ();
 sg13g2_fill_8 FILLER_0_91_144 ();
 sg13g2_fill_8 FILLER_0_91_152 ();
 sg13g2_fill_8 FILLER_0_91_160 ();
 sg13g2_fill_8 FILLER_0_91_168 ();
 sg13g2_fill_8 FILLER_0_91_176 ();
 sg13g2_fill_8 FILLER_0_91_184 ();
 sg13g2_fill_8 FILLER_0_91_192 ();
 sg13g2_fill_8 FILLER_0_91_200 ();
 sg13g2_fill_8 FILLER_0_91_208 ();
 sg13g2_fill_8 FILLER_0_91_216 ();
 sg13g2_fill_8 FILLER_0_91_224 ();
 sg13g2_fill_8 FILLER_0_91_232 ();
 sg13g2_fill_8 FILLER_0_91_240 ();
 sg13g2_fill_8 FILLER_0_91_248 ();
 sg13g2_fill_8 FILLER_0_91_256 ();
 sg13g2_fill_4 FILLER_0_91_264 ();
 sg13g2_fill_1 FILLER_0_91_268 ();
 sg13g2_fill_2 FILLER_0_91_295 ();
 sg13g2_fill_8 FILLER_0_91_318 ();
 sg13g2_fill_8 FILLER_0_91_326 ();
 sg13g2_fill_2 FILLER_0_91_334 ();
 sg13g2_fill_4 FILLER_0_91_341 ();
 sg13g2_fill_2 FILLER_0_91_345 ();
 sg13g2_fill_1 FILLER_0_91_347 ();
 sg13g2_fill_8 FILLER_0_91_352 ();
 sg13g2_fill_2 FILLER_0_91_360 ();
 sg13g2_fill_1 FILLER_0_91_362 ();
 sg13g2_fill_2 FILLER_0_91_369 ();
 sg13g2_fill_8 FILLER_0_91_376 ();
 sg13g2_fill_2 FILLER_0_91_410 ();
 sg13g2_fill_4 FILLER_0_91_417 ();
 sg13g2_fill_1 FILLER_0_91_421 ();
 sg13g2_fill_8 FILLER_0_91_427 ();
 sg13g2_fill_4 FILLER_0_91_435 ();
 sg13g2_fill_1 FILLER_0_91_439 ();
 sg13g2_fill_8 FILLER_0_91_445 ();
 sg13g2_fill_8 FILLER_0_91_453 ();
 sg13g2_fill_8 FILLER_0_91_461 ();
 sg13g2_fill_2 FILLER_0_91_469 ();
 sg13g2_fill_2 FILLER_0_91_497 ();
 sg13g2_fill_1 FILLER_0_91_499 ();
 sg13g2_fill_2 FILLER_0_91_505 ();
 sg13g2_fill_4 FILLER_0_91_513 ();
 sg13g2_fill_2 FILLER_0_91_517 ();
 sg13g2_fill_8 FILLER_0_91_545 ();
 sg13g2_fill_8 FILLER_0_91_553 ();
 sg13g2_fill_4 FILLER_0_91_561 ();
 sg13g2_fill_8 FILLER_0_91_570 ();
 sg13g2_fill_8 FILLER_0_91_578 ();
 sg13g2_fill_4 FILLER_0_91_586 ();
 sg13g2_fill_8 FILLER_0_91_595 ();
 sg13g2_fill_2 FILLER_0_91_629 ();
 sg13g2_fill_8 FILLER_0_91_657 ();
 sg13g2_fill_2 FILLER_0_91_665 ();
 sg13g2_fill_8 FILLER_0_91_672 ();
 sg13g2_fill_4 FILLER_0_91_680 ();
 sg13g2_fill_2 FILLER_0_91_684 ();
 sg13g2_fill_2 FILLER_0_91_691 ();
 sg13g2_fill_2 FILLER_0_91_698 ();
 sg13g2_fill_8 FILLER_0_91_705 ();
 sg13g2_fill_8 FILLER_0_91_713 ();
 sg13g2_fill_2 FILLER_0_91_726 ();
 sg13g2_fill_4 FILLER_0_91_733 ();
 sg13g2_fill_1 FILLER_0_91_737 ();
 sg13g2_fill_2 FILLER_0_91_743 ();
 sg13g2_fill_8 FILLER_0_91_771 ();
 sg13g2_fill_8 FILLER_0_91_789 ();
 sg13g2_fill_8 FILLER_0_91_797 ();
 sg13g2_fill_8 FILLER_0_91_805 ();
 sg13g2_fill_4 FILLER_0_91_813 ();
 sg13g2_fill_2 FILLER_0_91_821 ();
 sg13g2_fill_8 FILLER_0_91_827 ();
 sg13g2_fill_8 FILLER_0_91_835 ();
 sg13g2_fill_1 FILLER_0_91_843 ();
 sg13g2_fill_8 FILLER_0_91_852 ();
 sg13g2_fill_4 FILLER_0_91_860 ();
 sg13g2_fill_2 FILLER_0_91_864 ();
 sg13g2_fill_2 FILLER_0_91_871 ();
 sg13g2_fill_8 FILLER_0_91_876 ();
 sg13g2_fill_8 FILLER_0_91_884 ();
 sg13g2_fill_8 FILLER_0_91_892 ();
 sg13g2_fill_1 FILLER_0_91_900 ();
 sg13g2_fill_2 FILLER_0_91_904 ();
 sg13g2_fill_1 FILLER_0_91_906 ();
 sg13g2_fill_4 FILLER_0_91_912 ();
 sg13g2_fill_1 FILLER_0_91_916 ();
 sg13g2_fill_4 FILLER_0_91_927 ();
 sg13g2_fill_2 FILLER_0_91_931 ();
 sg13g2_fill_2 FILLER_0_91_943 ();
 sg13g2_fill_2 FILLER_0_91_950 ();
 sg13g2_fill_1 FILLER_0_91_952 ();
 sg13g2_fill_8 FILLER_0_91_963 ();
 sg13g2_fill_8 FILLER_0_91_971 ();
 sg13g2_fill_4 FILLER_0_91_979 ();
 sg13g2_fill_2 FILLER_0_91_983 ();
 sg13g2_fill_1 FILLER_0_91_985 ();
 sg13g2_fill_8 FILLER_0_91_991 ();
 sg13g2_fill_4 FILLER_0_91_999 ();
 sg13g2_fill_2 FILLER_0_91_1003 ();
 sg13g2_fill_1 FILLER_0_91_1005 ();
 sg13g2_fill_8 FILLER_0_91_1012 ();
 sg13g2_fill_8 FILLER_0_91_1020 ();
 sg13g2_fill_4 FILLER_0_91_1028 ();
 sg13g2_fill_1 FILLER_0_91_1032 ();
 sg13g2_fill_2 FILLER_0_91_1038 ();
 sg13g2_fill_8 FILLER_0_91_1045 ();
 sg13g2_fill_8 FILLER_0_91_1053 ();
 sg13g2_fill_2 FILLER_0_91_1061 ();
 sg13g2_fill_1 FILLER_0_91_1063 ();
 sg13g2_fill_8 FILLER_0_91_1068 ();
 sg13g2_fill_8 FILLER_0_91_1076 ();
 sg13g2_fill_2 FILLER_0_91_1084 ();
 sg13g2_fill_1 FILLER_0_91_1086 ();
 sg13g2_fill_2 FILLER_0_91_1092 ();
 sg13g2_fill_8 FILLER_0_91_1102 ();
 sg13g2_fill_8 FILLER_0_91_1110 ();
 sg13g2_fill_8 FILLER_0_91_1118 ();
 sg13g2_fill_8 FILLER_0_91_1126 ();
 sg13g2_fill_8 FILLER_0_91_1134 ();
 sg13g2_fill_8 FILLER_0_91_1142 ();
 sg13g2_fill_8 FILLER_0_91_1150 ();
 sg13g2_fill_8 FILLER_0_91_1158 ();
 sg13g2_fill_2 FILLER_0_91_1166 ();
 sg13g2_fill_1 FILLER_0_91_1168 ();
 sg13g2_fill_8 FILLER_0_91_1174 ();
 sg13g2_fill_4 FILLER_0_91_1182 ();
 sg13g2_fill_1 FILLER_0_91_1186 ();
 sg13g2_fill_8 FILLER_0_91_1195 ();
 sg13g2_fill_8 FILLER_0_91_1203 ();
 sg13g2_fill_8 FILLER_0_91_1211 ();
 sg13g2_fill_1 FILLER_0_91_1219 ();
 sg13g2_fill_4 FILLER_0_91_1224 ();
 sg13g2_fill_2 FILLER_0_91_1228 ();
 sg13g2_fill_1 FILLER_0_91_1230 ();
 sg13g2_fill_8 FILLER_0_91_1235 ();
 sg13g2_fill_2 FILLER_0_91_1247 ();
 sg13g2_fill_4 FILLER_0_91_1253 ();
 sg13g2_fill_1 FILLER_0_91_1257 ();
 sg13g2_fill_2 FILLER_0_91_1262 ();
 sg13g2_fill_2 FILLER_0_91_1270 ();
 sg13g2_fill_8 FILLER_0_91_1277 ();
 sg13g2_fill_8 FILLER_0_91_1289 ();
 sg13g2_fill_8 FILLER_0_92_0 ();
 sg13g2_fill_8 FILLER_0_92_8 ();
 sg13g2_fill_8 FILLER_0_92_16 ();
 sg13g2_fill_8 FILLER_0_92_24 ();
 sg13g2_fill_8 FILLER_0_92_32 ();
 sg13g2_fill_8 FILLER_0_92_40 ();
 sg13g2_fill_8 FILLER_0_92_48 ();
 sg13g2_fill_8 FILLER_0_92_56 ();
 sg13g2_fill_8 FILLER_0_92_64 ();
 sg13g2_fill_8 FILLER_0_92_72 ();
 sg13g2_fill_8 FILLER_0_92_80 ();
 sg13g2_fill_8 FILLER_0_92_88 ();
 sg13g2_fill_8 FILLER_0_92_96 ();
 sg13g2_fill_8 FILLER_0_92_104 ();
 sg13g2_fill_8 FILLER_0_92_112 ();
 sg13g2_fill_8 FILLER_0_92_120 ();
 sg13g2_fill_8 FILLER_0_92_128 ();
 sg13g2_fill_8 FILLER_0_92_136 ();
 sg13g2_fill_8 FILLER_0_92_144 ();
 sg13g2_fill_8 FILLER_0_92_152 ();
 sg13g2_fill_8 FILLER_0_92_160 ();
 sg13g2_fill_8 FILLER_0_92_168 ();
 sg13g2_fill_8 FILLER_0_92_176 ();
 sg13g2_fill_8 FILLER_0_92_184 ();
 sg13g2_fill_8 FILLER_0_92_192 ();
 sg13g2_fill_8 FILLER_0_92_200 ();
 sg13g2_fill_8 FILLER_0_92_208 ();
 sg13g2_fill_8 FILLER_0_92_216 ();
 sg13g2_fill_8 FILLER_0_92_224 ();
 sg13g2_fill_8 FILLER_0_92_232 ();
 sg13g2_fill_8 FILLER_0_92_240 ();
 sg13g2_fill_4 FILLER_0_92_248 ();
 sg13g2_fill_2 FILLER_0_92_257 ();
 sg13g2_fill_2 FILLER_0_92_263 ();
 sg13g2_fill_2 FILLER_0_92_269 ();
 sg13g2_fill_2 FILLER_0_92_297 ();
 sg13g2_fill_2 FILLER_0_92_325 ();
 sg13g2_fill_8 FILLER_0_92_332 ();
 sg13g2_fill_8 FILLER_0_92_340 ();
 sg13g2_fill_8 FILLER_0_92_353 ();
 sg13g2_fill_1 FILLER_0_92_361 ();
 sg13g2_fill_2 FILLER_0_92_367 ();
 sg13g2_fill_8 FILLER_0_92_374 ();
 sg13g2_fill_8 FILLER_0_92_382 ();
 sg13g2_fill_8 FILLER_0_92_390 ();
 sg13g2_fill_8 FILLER_0_92_398 ();
 sg13g2_fill_1 FILLER_0_92_406 ();
 sg13g2_fill_4 FILLER_0_92_412 ();
 sg13g2_fill_2 FILLER_0_92_416 ();
 sg13g2_fill_1 FILLER_0_92_418 ();
 sg13g2_fill_8 FILLER_0_92_445 ();
 sg13g2_fill_4 FILLER_0_92_453 ();
 sg13g2_fill_2 FILLER_0_92_457 ();
 sg13g2_fill_1 FILLER_0_92_459 ();
 sg13g2_fill_8 FILLER_0_92_465 ();
 sg13g2_fill_8 FILLER_0_92_477 ();
 sg13g2_fill_8 FILLER_0_92_485 ();
 sg13g2_fill_2 FILLER_0_92_493 ();
 sg13g2_fill_8 FILLER_0_92_500 ();
 sg13g2_fill_8 FILLER_0_92_508 ();
 sg13g2_fill_8 FILLER_0_92_516 ();
 sg13g2_fill_8 FILLER_0_92_524 ();
 sg13g2_fill_8 FILLER_0_92_532 ();
 sg13g2_fill_8 FILLER_0_92_540 ();
 sg13g2_fill_8 FILLER_0_92_548 ();
 sg13g2_fill_8 FILLER_0_92_556 ();
 sg13g2_fill_8 FILLER_0_92_564 ();
 sg13g2_fill_4 FILLER_0_92_572 ();
 sg13g2_fill_8 FILLER_0_92_583 ();
 sg13g2_fill_4 FILLER_0_92_591 ();
 sg13g2_fill_2 FILLER_0_92_595 ();
 sg13g2_fill_2 FILLER_0_92_602 ();
 sg13g2_fill_2 FILLER_0_92_608 ();
 sg13g2_fill_2 FILLER_0_92_615 ();
 sg13g2_fill_2 FILLER_0_92_627 ();
 sg13g2_fill_8 FILLER_0_92_634 ();
 sg13g2_fill_8 FILLER_0_92_652 ();
 sg13g2_fill_4 FILLER_0_92_660 ();
 sg13g2_fill_2 FILLER_0_92_664 ();
 sg13g2_fill_1 FILLER_0_92_666 ();
 sg13g2_fill_2 FILLER_0_92_672 ();
 sg13g2_fill_1 FILLER_0_92_674 ();
 sg13g2_fill_8 FILLER_0_92_683 ();
 sg13g2_fill_8 FILLER_0_92_691 ();
 sg13g2_fill_4 FILLER_0_92_699 ();
 sg13g2_fill_2 FILLER_0_92_703 ();
 sg13g2_fill_4 FILLER_0_92_715 ();
 sg13g2_fill_2 FILLER_0_92_719 ();
 sg13g2_fill_4 FILLER_0_92_725 ();
 sg13g2_fill_1 FILLER_0_92_729 ();
 sg13g2_fill_2 FILLER_0_92_756 ();
 sg13g2_fill_2 FILLER_0_92_764 ();
 sg13g2_fill_1 FILLER_0_92_766 ();
 sg13g2_fill_2 FILLER_0_92_773 ();
 sg13g2_fill_1 FILLER_0_92_775 ();
 sg13g2_fill_2 FILLER_0_92_781 ();
 sg13g2_fill_1 FILLER_0_92_783 ();
 sg13g2_fill_2 FILLER_0_92_810 ();
 sg13g2_fill_2 FILLER_0_92_816 ();
 sg13g2_fill_1 FILLER_0_92_818 ();
 sg13g2_fill_2 FILLER_0_92_825 ();
 sg13g2_fill_8 FILLER_0_92_832 ();
 sg13g2_fill_1 FILLER_0_92_840 ();
 sg13g2_fill_4 FILLER_0_92_846 ();
 sg13g2_fill_1 FILLER_0_92_850 ();
 sg13g2_fill_8 FILLER_0_92_856 ();
 sg13g2_fill_2 FILLER_0_92_873 ();
 sg13g2_fill_2 FILLER_0_92_880 ();
 sg13g2_fill_8 FILLER_0_92_891 ();
 sg13g2_fill_8 FILLER_0_92_899 ();
 sg13g2_fill_8 FILLER_0_92_907 ();
 sg13g2_fill_4 FILLER_0_92_915 ();
 sg13g2_fill_1 FILLER_0_92_919 ();
 sg13g2_fill_8 FILLER_0_92_930 ();
 sg13g2_fill_1 FILLER_0_92_938 ();
 sg13g2_fill_8 FILLER_0_92_943 ();
 sg13g2_fill_2 FILLER_0_92_951 ();
 sg13g2_fill_8 FILLER_0_92_957 ();
 sg13g2_fill_2 FILLER_0_92_965 ();
 sg13g2_fill_1 FILLER_0_92_967 ();
 sg13g2_fill_4 FILLER_0_92_978 ();
 sg13g2_fill_2 FILLER_0_92_982 ();
 sg13g2_fill_1 FILLER_0_92_984 ();
 sg13g2_fill_8 FILLER_0_92_989 ();
 sg13g2_fill_8 FILLER_0_92_997 ();
 sg13g2_fill_4 FILLER_0_92_1005 ();
 sg13g2_fill_4 FILLER_0_92_1014 ();
 sg13g2_fill_2 FILLER_0_92_1018 ();
 sg13g2_fill_1 FILLER_0_92_1020 ();
 sg13g2_fill_8 FILLER_0_92_1025 ();
 sg13g2_fill_1 FILLER_0_92_1033 ();
 sg13g2_fill_8 FILLER_0_92_1040 ();
 sg13g2_fill_8 FILLER_0_92_1048 ();
 sg13g2_fill_8 FILLER_0_92_1056 ();
 sg13g2_fill_2 FILLER_0_92_1064 ();
 sg13g2_fill_8 FILLER_0_92_1071 ();
 sg13g2_fill_8 FILLER_0_92_1079 ();
 sg13g2_fill_8 FILLER_0_92_1087 ();
 sg13g2_fill_8 FILLER_0_92_1095 ();
 sg13g2_fill_8 FILLER_0_92_1103 ();
 sg13g2_fill_8 FILLER_0_92_1111 ();
 sg13g2_fill_8 FILLER_0_92_1119 ();
 sg13g2_fill_8 FILLER_0_92_1127 ();
 sg13g2_fill_4 FILLER_0_92_1135 ();
 sg13g2_fill_8 FILLER_0_92_1144 ();
 sg13g2_fill_8 FILLER_0_92_1152 ();
 sg13g2_fill_2 FILLER_0_92_1165 ();
 sg13g2_fill_2 FILLER_0_92_1171 ();
 sg13g2_fill_2 FILLER_0_92_1178 ();
 sg13g2_fill_8 FILLER_0_92_1184 ();
 sg13g2_fill_4 FILLER_0_92_1197 ();
 sg13g2_fill_8 FILLER_0_92_1209 ();
 sg13g2_fill_8 FILLER_0_92_1217 ();
 sg13g2_fill_8 FILLER_0_92_1225 ();
 sg13g2_fill_8 FILLER_0_92_1233 ();
 sg13g2_fill_4 FILLER_0_92_1241 ();
 sg13g2_fill_2 FILLER_0_92_1245 ();
 sg13g2_fill_2 FILLER_0_92_1253 ();
 sg13g2_fill_8 FILLER_0_92_1259 ();
 sg13g2_fill_2 FILLER_0_92_1272 ();
 sg13g2_fill_2 FILLER_0_92_1278 ();
 sg13g2_fill_2 FILLER_0_92_1284 ();
 sg13g2_fill_2 FILLER_0_92_1290 ();
 sg13g2_fill_1 FILLER_0_92_1296 ();
 sg13g2_fill_8 FILLER_0_93_0 ();
 sg13g2_fill_8 FILLER_0_93_8 ();
 sg13g2_fill_8 FILLER_0_93_16 ();
 sg13g2_fill_8 FILLER_0_93_24 ();
 sg13g2_fill_8 FILLER_0_93_32 ();
 sg13g2_fill_8 FILLER_0_93_40 ();
 sg13g2_fill_8 FILLER_0_93_48 ();
 sg13g2_fill_8 FILLER_0_93_56 ();
 sg13g2_fill_8 FILLER_0_93_64 ();
 sg13g2_fill_8 FILLER_0_93_72 ();
 sg13g2_fill_8 FILLER_0_93_80 ();
 sg13g2_fill_8 FILLER_0_93_88 ();
 sg13g2_fill_8 FILLER_0_93_96 ();
 sg13g2_fill_8 FILLER_0_93_104 ();
 sg13g2_fill_8 FILLER_0_93_112 ();
 sg13g2_fill_8 FILLER_0_93_120 ();
 sg13g2_fill_8 FILLER_0_93_128 ();
 sg13g2_fill_8 FILLER_0_93_136 ();
 sg13g2_fill_8 FILLER_0_93_144 ();
 sg13g2_fill_8 FILLER_0_93_152 ();
 sg13g2_fill_8 FILLER_0_93_160 ();
 sg13g2_fill_8 FILLER_0_93_168 ();
 sg13g2_fill_8 FILLER_0_93_176 ();
 sg13g2_fill_8 FILLER_0_93_184 ();
 sg13g2_fill_8 FILLER_0_93_192 ();
 sg13g2_fill_8 FILLER_0_93_200 ();
 sg13g2_fill_8 FILLER_0_93_208 ();
 sg13g2_fill_8 FILLER_0_93_216 ();
 sg13g2_fill_8 FILLER_0_93_224 ();
 sg13g2_fill_8 FILLER_0_93_232 ();
 sg13g2_fill_8 FILLER_0_93_240 ();
 sg13g2_fill_2 FILLER_0_93_248 ();
 sg13g2_fill_1 FILLER_0_93_250 ();
 sg13g2_fill_4 FILLER_0_93_277 ();
 sg13g2_fill_2 FILLER_0_93_286 ();
 sg13g2_fill_1 FILLER_0_93_288 ();
 sg13g2_fill_2 FILLER_0_93_293 ();
 sg13g2_fill_8 FILLER_0_93_316 ();
 sg13g2_fill_4 FILLER_0_93_324 ();
 sg13g2_fill_8 FILLER_0_93_332 ();
 sg13g2_fill_1 FILLER_0_93_340 ();
 sg13g2_fill_2 FILLER_0_93_367 ();
 sg13g2_fill_1 FILLER_0_93_369 ();
 sg13g2_fill_8 FILLER_0_93_374 ();
 sg13g2_fill_8 FILLER_0_93_382 ();
 sg13g2_fill_8 FILLER_0_93_390 ();
 sg13g2_fill_2 FILLER_0_93_398 ();
 sg13g2_fill_1 FILLER_0_93_400 ();
 sg13g2_fill_8 FILLER_0_93_405 ();
 sg13g2_fill_8 FILLER_0_93_413 ();
 sg13g2_fill_8 FILLER_0_93_421 ();
 sg13g2_fill_8 FILLER_0_93_429 ();
 sg13g2_fill_8 FILLER_0_93_437 ();
 sg13g2_fill_8 FILLER_0_93_445 ();
 sg13g2_fill_4 FILLER_0_93_479 ();
 sg13g2_fill_2 FILLER_0_93_483 ();
 sg13g2_fill_1 FILLER_0_93_485 ();
 sg13g2_fill_4 FILLER_0_93_491 ();
 sg13g2_fill_2 FILLER_0_93_495 ();
 sg13g2_fill_2 FILLER_0_93_503 ();
 sg13g2_fill_8 FILLER_0_93_512 ();
 sg13g2_fill_8 FILLER_0_93_520 ();
 sg13g2_fill_8 FILLER_0_93_528 ();
 sg13g2_fill_8 FILLER_0_93_536 ();
 sg13g2_fill_8 FILLER_0_93_544 ();
 sg13g2_fill_8 FILLER_0_93_552 ();
 sg13g2_fill_4 FILLER_0_93_560 ();
 sg13g2_fill_2 FILLER_0_93_564 ();
 sg13g2_fill_8 FILLER_0_93_578 ();
 sg13g2_fill_8 FILLER_0_93_586 ();
 sg13g2_fill_8 FILLER_0_93_594 ();
 sg13g2_fill_2 FILLER_0_93_607 ();
 sg13g2_fill_4 FILLER_0_93_613 ();
 sg13g2_fill_2 FILLER_0_93_617 ();
 sg13g2_fill_1 FILLER_0_93_619 ();
 sg13g2_fill_2 FILLER_0_93_626 ();
 sg13g2_fill_8 FILLER_0_93_633 ();
 sg13g2_fill_8 FILLER_0_93_641 ();
 sg13g2_fill_8 FILLER_0_93_649 ();
 sg13g2_fill_8 FILLER_0_93_657 ();
 sg13g2_fill_4 FILLER_0_93_665 ();
 sg13g2_fill_1 FILLER_0_93_669 ();
 sg13g2_fill_4 FILLER_0_93_680 ();
 sg13g2_fill_2 FILLER_0_93_684 ();
 sg13g2_fill_4 FILLER_0_93_690 ();
 sg13g2_fill_8 FILLER_0_93_698 ();
 sg13g2_fill_8 FILLER_0_93_706 ();
 sg13g2_fill_4 FILLER_0_93_714 ();
 sg13g2_fill_1 FILLER_0_93_718 ();
 sg13g2_fill_8 FILLER_0_93_729 ();
 sg13g2_fill_4 FILLER_0_93_737 ();
 sg13g2_fill_2 FILLER_0_93_741 ();
 sg13g2_fill_1 FILLER_0_93_743 ();
 sg13g2_fill_4 FILLER_0_93_754 ();
 sg13g2_fill_1 FILLER_0_93_758 ();
 sg13g2_fill_4 FILLER_0_93_769 ();
 sg13g2_fill_1 FILLER_0_93_773 ();
 sg13g2_fill_8 FILLER_0_93_780 ();
 sg13g2_fill_8 FILLER_0_93_788 ();
 sg13g2_fill_2 FILLER_0_93_802 ();
 sg13g2_fill_4 FILLER_0_93_808 ();
 sg13g2_fill_4 FILLER_0_93_816 ();
 sg13g2_fill_1 FILLER_0_93_820 ();
 sg13g2_fill_2 FILLER_0_93_825 ();
 sg13g2_fill_2 FILLER_0_93_831 ();
 sg13g2_fill_2 FILLER_0_93_837 ();
 sg13g2_fill_1 FILLER_0_93_839 ();
 sg13g2_fill_8 FILLER_0_93_844 ();
 sg13g2_fill_8 FILLER_0_93_852 ();
 sg13g2_fill_4 FILLER_0_93_860 ();
 sg13g2_fill_2 FILLER_0_93_864 ();
 sg13g2_fill_2 FILLER_0_93_873 ();
 sg13g2_fill_4 FILLER_0_93_880 ();
 sg13g2_fill_2 FILLER_0_93_884 ();
 sg13g2_fill_8 FILLER_0_93_891 ();
 sg13g2_fill_8 FILLER_0_93_899 ();
 sg13g2_fill_8 FILLER_0_93_907 ();
 sg13g2_fill_8 FILLER_0_93_915 ();
 sg13g2_fill_8 FILLER_0_93_933 ();
 sg13g2_fill_4 FILLER_0_93_946 ();
 sg13g2_fill_2 FILLER_0_93_955 ();
 sg13g2_fill_2 FILLER_0_93_961 ();
 sg13g2_fill_1 FILLER_0_93_963 ();
 sg13g2_fill_2 FILLER_0_93_968 ();
 sg13g2_fill_8 FILLER_0_93_974 ();
 sg13g2_fill_1 FILLER_0_93_982 ();
 sg13g2_fill_4 FILLER_0_93_988 ();
 sg13g2_fill_2 FILLER_0_93_992 ();
 sg13g2_fill_1 FILLER_0_93_994 ();
 sg13g2_fill_2 FILLER_0_93_1000 ();
 sg13g2_fill_2 FILLER_0_93_1012 ();
 sg13g2_fill_2 FILLER_0_93_1020 ();
 sg13g2_fill_1 FILLER_0_93_1022 ();
 sg13g2_fill_4 FILLER_0_93_1027 ();
 sg13g2_fill_2 FILLER_0_93_1031 ();
 sg13g2_fill_1 FILLER_0_93_1033 ();
 sg13g2_fill_2 FILLER_0_93_1039 ();
 sg13g2_fill_2 FILLER_0_93_1047 ();
 sg13g2_fill_4 FILLER_0_93_1055 ();
 sg13g2_fill_2 FILLER_0_93_1059 ();
 sg13g2_fill_1 FILLER_0_93_1061 ();
 sg13g2_fill_4 FILLER_0_93_1070 ();
 sg13g2_fill_8 FILLER_0_93_1081 ();
 sg13g2_fill_8 FILLER_0_93_1089 ();
 sg13g2_fill_8 FILLER_0_93_1097 ();
 sg13g2_fill_8 FILLER_0_93_1105 ();
 sg13g2_fill_4 FILLER_0_93_1113 ();
 sg13g2_fill_1 FILLER_0_93_1117 ();
 sg13g2_fill_2 FILLER_0_93_1122 ();
 sg13g2_fill_1 FILLER_0_93_1124 ();
 sg13g2_fill_4 FILLER_0_93_1129 ();
 sg13g2_fill_4 FILLER_0_93_1138 ();
 sg13g2_fill_4 FILLER_0_93_1150 ();
 sg13g2_fill_2 FILLER_0_93_1159 ();
 sg13g2_fill_1 FILLER_0_93_1161 ();
 sg13g2_fill_2 FILLER_0_93_1166 ();
 sg13g2_fill_2 FILLER_0_93_1173 ();
 sg13g2_fill_4 FILLER_0_93_1178 ();
 sg13g2_fill_1 FILLER_0_93_1182 ();
 sg13g2_fill_2 FILLER_0_93_1188 ();
 sg13g2_fill_2 FILLER_0_93_1197 ();
 sg13g2_fill_4 FILLER_0_93_1209 ();
 sg13g2_fill_1 FILLER_0_93_1213 ();
 sg13g2_fill_8 FILLER_0_93_1221 ();
 sg13g2_fill_2 FILLER_0_93_1229 ();
 sg13g2_fill_1 FILLER_0_93_1231 ();
 sg13g2_fill_2 FILLER_0_93_1240 ();
 sg13g2_fill_1 FILLER_0_93_1242 ();
 sg13g2_fill_2 FILLER_0_93_1251 ();
 sg13g2_fill_4 FILLER_0_93_1260 ();
 sg13g2_fill_2 FILLER_0_93_1268 ();
 sg13g2_fill_4 FILLER_0_93_1275 ();
 sg13g2_fill_2 FILLER_0_93_1279 ();
 sg13g2_fill_8 FILLER_0_93_1286 ();
 sg13g2_fill_2 FILLER_0_93_1294 ();
 sg13g2_fill_1 FILLER_0_93_1296 ();
 sg13g2_fill_8 FILLER_0_94_0 ();
 sg13g2_fill_8 FILLER_0_94_8 ();
 sg13g2_fill_8 FILLER_0_94_16 ();
 sg13g2_fill_8 FILLER_0_94_24 ();
 sg13g2_fill_8 FILLER_0_94_32 ();
 sg13g2_fill_8 FILLER_0_94_40 ();
 sg13g2_fill_8 FILLER_0_94_48 ();
 sg13g2_fill_8 FILLER_0_94_56 ();
 sg13g2_fill_8 FILLER_0_94_64 ();
 sg13g2_fill_8 FILLER_0_94_72 ();
 sg13g2_fill_8 FILLER_0_94_80 ();
 sg13g2_fill_8 FILLER_0_94_88 ();
 sg13g2_fill_8 FILLER_0_94_96 ();
 sg13g2_fill_8 FILLER_0_94_104 ();
 sg13g2_fill_8 FILLER_0_94_112 ();
 sg13g2_fill_8 FILLER_0_94_120 ();
 sg13g2_fill_8 FILLER_0_94_128 ();
 sg13g2_fill_8 FILLER_0_94_136 ();
 sg13g2_fill_8 FILLER_0_94_144 ();
 sg13g2_fill_8 FILLER_0_94_152 ();
 sg13g2_fill_8 FILLER_0_94_160 ();
 sg13g2_fill_8 FILLER_0_94_168 ();
 sg13g2_fill_8 FILLER_0_94_176 ();
 sg13g2_fill_8 FILLER_0_94_184 ();
 sg13g2_fill_8 FILLER_0_94_192 ();
 sg13g2_fill_8 FILLER_0_94_200 ();
 sg13g2_fill_8 FILLER_0_94_208 ();
 sg13g2_fill_8 FILLER_0_94_216 ();
 sg13g2_fill_8 FILLER_0_94_224 ();
 sg13g2_fill_8 FILLER_0_94_232 ();
 sg13g2_fill_8 FILLER_0_94_240 ();
 sg13g2_fill_8 FILLER_0_94_248 ();
 sg13g2_fill_8 FILLER_0_94_256 ();
 sg13g2_fill_8 FILLER_0_94_264 ();
 sg13g2_fill_8 FILLER_0_94_272 ();
 sg13g2_fill_8 FILLER_0_94_280 ();
 sg13g2_fill_8 FILLER_0_94_288 ();
 sg13g2_fill_8 FILLER_0_94_296 ();
 sg13g2_fill_8 FILLER_0_94_304 ();
 sg13g2_fill_8 FILLER_0_94_312 ();
 sg13g2_fill_8 FILLER_0_94_320 ();
 sg13g2_fill_2 FILLER_0_94_328 ();
 sg13g2_fill_1 FILLER_0_94_330 ();
 sg13g2_fill_4 FILLER_0_94_336 ();
 sg13g2_fill_2 FILLER_0_94_340 ();
 sg13g2_fill_8 FILLER_0_94_346 ();
 sg13g2_fill_8 FILLER_0_94_354 ();
 sg13g2_fill_8 FILLER_0_94_362 ();
 sg13g2_fill_8 FILLER_0_94_370 ();
 sg13g2_fill_4 FILLER_0_94_378 ();
 sg13g2_fill_1 FILLER_0_94_382 ();
 sg13g2_fill_2 FILLER_0_94_388 ();
 sg13g2_fill_4 FILLER_0_94_416 ();
 sg13g2_fill_1 FILLER_0_94_420 ();
 sg13g2_fill_2 FILLER_0_94_425 ();
 sg13g2_fill_8 FILLER_0_94_437 ();
 sg13g2_fill_8 FILLER_0_94_445 ();
 sg13g2_fill_8 FILLER_0_94_453 ();
 sg13g2_fill_4 FILLER_0_94_461 ();
 sg13g2_fill_1 FILLER_0_94_465 ();
 sg13g2_fill_2 FILLER_0_94_471 ();
 sg13g2_fill_2 FILLER_0_94_479 ();
 sg13g2_fill_8 FILLER_0_94_485 ();
 sg13g2_fill_8 FILLER_0_94_493 ();
 sg13g2_fill_4 FILLER_0_94_501 ();
 sg13g2_fill_1 FILLER_0_94_505 ();
 sg13g2_fill_8 FILLER_0_94_511 ();
 sg13g2_fill_8 FILLER_0_94_519 ();
 sg13g2_fill_4 FILLER_0_94_531 ();
 sg13g2_fill_2 FILLER_0_94_541 ();
 sg13g2_fill_8 FILLER_0_94_548 ();
 sg13g2_fill_4 FILLER_0_94_556 ();
 sg13g2_fill_2 FILLER_0_94_560 ();
 sg13g2_fill_8 FILLER_0_94_567 ();
 sg13g2_fill_8 FILLER_0_94_575 ();
 sg13g2_fill_8 FILLER_0_94_583 ();
 sg13g2_fill_8 FILLER_0_94_591 ();
 sg13g2_fill_4 FILLER_0_94_599 ();
 sg13g2_fill_8 FILLER_0_94_608 ();
 sg13g2_fill_8 FILLER_0_94_616 ();
 sg13g2_fill_8 FILLER_0_94_624 ();
 sg13g2_fill_8 FILLER_0_94_632 ();
 sg13g2_fill_8 FILLER_0_94_640 ();
 sg13g2_fill_2 FILLER_0_94_648 ();
 sg13g2_fill_1 FILLER_0_94_650 ();
 sg13g2_fill_8 FILLER_0_94_661 ();
 sg13g2_fill_1 FILLER_0_94_669 ();
 sg13g2_fill_2 FILLER_0_94_696 ();
 sg13g2_fill_8 FILLER_0_94_724 ();
 sg13g2_fill_8 FILLER_0_94_732 ();
 sg13g2_fill_4 FILLER_0_94_740 ();
 sg13g2_fill_2 FILLER_0_94_744 ();
 sg13g2_fill_2 FILLER_0_94_751 ();
 sg13g2_fill_2 FILLER_0_94_757 ();
 sg13g2_fill_4 FILLER_0_94_769 ();
 sg13g2_fill_1 FILLER_0_94_773 ();
 sg13g2_fill_4 FILLER_0_94_780 ();
 sg13g2_fill_2 FILLER_0_94_794 ();
 sg13g2_fill_2 FILLER_0_94_801 ();
 sg13g2_fill_1 FILLER_0_94_803 ();
 sg13g2_fill_2 FILLER_0_94_809 ();
 sg13g2_fill_1 FILLER_0_94_811 ();
 sg13g2_fill_2 FILLER_0_94_816 ();
 sg13g2_fill_2 FILLER_0_94_822 ();
 sg13g2_fill_2 FILLER_0_94_828 ();
 sg13g2_fill_8 FILLER_0_94_834 ();
 sg13g2_fill_4 FILLER_0_94_842 ();
 sg13g2_fill_2 FILLER_0_94_846 ();
 sg13g2_fill_8 FILLER_0_94_852 ();
 sg13g2_fill_8 FILLER_0_94_860 ();
 sg13g2_fill_8 FILLER_0_94_868 ();
 sg13g2_fill_2 FILLER_0_94_876 ();
 sg13g2_fill_2 FILLER_0_94_883 ();
 sg13g2_fill_8 FILLER_0_94_890 ();
 sg13g2_fill_8 FILLER_0_94_898 ();
 sg13g2_fill_8 FILLER_0_94_906 ();
 sg13g2_fill_4 FILLER_0_94_914 ();
 sg13g2_fill_1 FILLER_0_94_918 ();
 sg13g2_fill_8 FILLER_0_94_929 ();
 sg13g2_fill_4 FILLER_0_94_937 ();
 sg13g2_fill_4 FILLER_0_94_946 ();
 sg13g2_fill_2 FILLER_0_94_950 ();
 sg13g2_fill_2 FILLER_0_94_957 ();
 sg13g2_fill_2 FILLER_0_94_964 ();
 sg13g2_fill_8 FILLER_0_94_971 ();
 sg13g2_fill_8 FILLER_0_94_979 ();
 sg13g2_fill_8 FILLER_0_94_987 ();
 sg13g2_fill_1 FILLER_0_94_995 ();
 sg13g2_fill_8 FILLER_0_94_1001 ();
 sg13g2_fill_8 FILLER_0_94_1009 ();
 sg13g2_fill_1 FILLER_0_94_1017 ();
 sg13g2_fill_4 FILLER_0_94_1022 ();
 sg13g2_fill_1 FILLER_0_94_1026 ();
 sg13g2_fill_4 FILLER_0_94_1032 ();
 sg13g2_fill_2 FILLER_0_94_1036 ();
 sg13g2_fill_1 FILLER_0_94_1038 ();
 sg13g2_fill_2 FILLER_0_94_1043 ();
 sg13g2_fill_4 FILLER_0_94_1049 ();
 sg13g2_fill_1 FILLER_0_94_1053 ();
 sg13g2_fill_4 FILLER_0_94_1058 ();
 sg13g2_fill_2 FILLER_0_94_1062 ();
 sg13g2_fill_2 FILLER_0_94_1068 ();
 sg13g2_fill_1 FILLER_0_94_1070 ();
 sg13g2_fill_4 FILLER_0_94_1076 ();
 sg13g2_fill_2 FILLER_0_94_1080 ();
 sg13g2_fill_8 FILLER_0_94_1087 ();
 sg13g2_fill_2 FILLER_0_94_1095 ();
 sg13g2_fill_4 FILLER_0_94_1102 ();
 sg13g2_fill_1 FILLER_0_94_1106 ();
 sg13g2_fill_4 FILLER_0_94_1115 ();
 sg13g2_fill_2 FILLER_0_94_1127 ();
 sg13g2_fill_2 FILLER_0_94_1132 ();
 sg13g2_fill_1 FILLER_0_94_1134 ();
 sg13g2_fill_8 FILLER_0_94_1139 ();
 sg13g2_fill_4 FILLER_0_94_1147 ();
 sg13g2_fill_2 FILLER_0_94_1151 ();
 sg13g2_fill_1 FILLER_0_94_1153 ();
 sg13g2_fill_4 FILLER_0_94_1158 ();
 sg13g2_fill_2 FILLER_0_94_1167 ();
 sg13g2_fill_2 FILLER_0_94_1174 ();
 sg13g2_fill_2 FILLER_0_94_1180 ();
 sg13g2_fill_4 FILLER_0_94_1186 ();
 sg13g2_fill_2 FILLER_0_94_1190 ();
 sg13g2_fill_1 FILLER_0_94_1192 ();
 sg13g2_fill_8 FILLER_0_94_1197 ();
 sg13g2_fill_8 FILLER_0_94_1205 ();
 sg13g2_fill_4 FILLER_0_94_1213 ();
 sg13g2_fill_1 FILLER_0_94_1217 ();
 sg13g2_fill_2 FILLER_0_94_1222 ();
 sg13g2_fill_2 FILLER_0_94_1229 ();
 sg13g2_fill_2 FILLER_0_94_1238 ();
 sg13g2_fill_4 FILLER_0_94_1245 ();
 sg13g2_fill_2 FILLER_0_94_1253 ();
 sg13g2_fill_2 FILLER_0_94_1259 ();
 sg13g2_fill_2 FILLER_0_94_1265 ();
 sg13g2_fill_2 FILLER_0_94_1272 ();
 sg13g2_fill_2 FILLER_0_94_1279 ();
 sg13g2_fill_2 FILLER_0_94_1286 ();
 sg13g2_fill_4 FILLER_0_94_1293 ();
 sg13g2_fill_8 FILLER_0_95_0 ();
 sg13g2_fill_8 FILLER_0_95_8 ();
 sg13g2_fill_8 FILLER_0_95_16 ();
 sg13g2_fill_8 FILLER_0_95_24 ();
 sg13g2_fill_8 FILLER_0_95_32 ();
 sg13g2_fill_8 FILLER_0_95_40 ();
 sg13g2_fill_8 FILLER_0_95_48 ();
 sg13g2_fill_8 FILLER_0_95_56 ();
 sg13g2_fill_8 FILLER_0_95_64 ();
 sg13g2_fill_8 FILLER_0_95_72 ();
 sg13g2_fill_8 FILLER_0_95_80 ();
 sg13g2_fill_8 FILLER_0_95_88 ();
 sg13g2_fill_8 FILLER_0_95_96 ();
 sg13g2_fill_8 FILLER_0_95_104 ();
 sg13g2_fill_8 FILLER_0_95_112 ();
 sg13g2_fill_8 FILLER_0_95_120 ();
 sg13g2_fill_8 FILLER_0_95_128 ();
 sg13g2_fill_8 FILLER_0_95_136 ();
 sg13g2_fill_8 FILLER_0_95_144 ();
 sg13g2_fill_8 FILLER_0_95_152 ();
 sg13g2_fill_8 FILLER_0_95_160 ();
 sg13g2_fill_8 FILLER_0_95_168 ();
 sg13g2_fill_8 FILLER_0_95_176 ();
 sg13g2_fill_8 FILLER_0_95_184 ();
 sg13g2_fill_8 FILLER_0_95_192 ();
 sg13g2_fill_8 FILLER_0_95_200 ();
 sg13g2_fill_8 FILLER_0_95_208 ();
 sg13g2_fill_8 FILLER_0_95_216 ();
 sg13g2_fill_8 FILLER_0_95_224 ();
 sg13g2_fill_8 FILLER_0_95_232 ();
 sg13g2_fill_1 FILLER_0_95_240 ();
 sg13g2_fill_4 FILLER_0_95_246 ();
 sg13g2_fill_8 FILLER_0_95_254 ();
 sg13g2_fill_8 FILLER_0_95_262 ();
 sg13g2_fill_8 FILLER_0_95_270 ();
 sg13g2_fill_2 FILLER_0_95_278 ();
 sg13g2_fill_8 FILLER_0_95_285 ();
 sg13g2_fill_8 FILLER_0_95_293 ();
 sg13g2_fill_8 FILLER_0_95_301 ();
 sg13g2_fill_8 FILLER_0_95_309 ();
 sg13g2_fill_8 FILLER_0_95_317 ();
 sg13g2_fill_1 FILLER_0_95_325 ();
 sg13g2_fill_8 FILLER_0_95_352 ();
 sg13g2_fill_8 FILLER_0_95_360 ();
 sg13g2_fill_4 FILLER_0_95_368 ();
 sg13g2_fill_1 FILLER_0_95_372 ();
 sg13g2_fill_2 FILLER_0_95_378 ();
 sg13g2_fill_8 FILLER_0_95_384 ();
 sg13g2_fill_8 FILLER_0_95_392 ();
 sg13g2_fill_8 FILLER_0_95_400 ();
 sg13g2_fill_4 FILLER_0_95_408 ();
 sg13g2_fill_1 FILLER_0_95_412 ();
 sg13g2_fill_2 FILLER_0_95_418 ();
 sg13g2_fill_4 FILLER_0_95_446 ();
 sg13g2_fill_2 FILLER_0_95_450 ();
 sg13g2_fill_1 FILLER_0_95_452 ();
 sg13g2_fill_4 FILLER_0_95_479 ();
 sg13g2_fill_1 FILLER_0_95_483 ();
 sg13g2_fill_4 FILLER_0_95_489 ();
 sg13g2_fill_2 FILLER_0_95_493 ();
 sg13g2_fill_8 FILLER_0_95_521 ();
 sg13g2_fill_1 FILLER_0_95_529 ();
 sg13g2_fill_8 FILLER_0_95_535 ();
 sg13g2_fill_8 FILLER_0_95_543 ();
 sg13g2_fill_8 FILLER_0_95_551 ();
 sg13g2_fill_2 FILLER_0_95_559 ();
 sg13g2_fill_1 FILLER_0_95_561 ();
 sg13g2_fill_2 FILLER_0_95_566 ();
 sg13g2_fill_4 FILLER_0_95_594 ();
 sg13g2_fill_2 FILLER_0_95_598 ();
 sg13g2_fill_1 FILLER_0_95_600 ();
 sg13g2_fill_8 FILLER_0_95_605 ();
 sg13g2_fill_8 FILLER_0_95_613 ();
 sg13g2_fill_2 FILLER_0_95_621 ();
 sg13g2_fill_8 FILLER_0_95_629 ();
 sg13g2_fill_4 FILLER_0_95_637 ();
 sg13g2_fill_4 FILLER_0_95_646 ();
 sg13g2_fill_2 FILLER_0_95_650 ();
 sg13g2_fill_2 FILLER_0_95_678 ();
 sg13g2_fill_8 FILLER_0_95_684 ();
 sg13g2_fill_2 FILLER_0_95_698 ();
 sg13g2_fill_2 FILLER_0_95_705 ();
 sg13g2_fill_2 FILLER_0_95_717 ();
 sg13g2_fill_8 FILLER_0_95_729 ();
 sg13g2_fill_8 FILLER_0_95_737 ();
 sg13g2_fill_8 FILLER_0_95_745 ();
 sg13g2_fill_8 FILLER_0_95_753 ();
 sg13g2_fill_4 FILLER_0_95_761 ();
 sg13g2_fill_2 FILLER_0_95_791 ();
 sg13g2_fill_4 FILLER_0_95_798 ();
 sg13g2_fill_2 FILLER_0_95_802 ();
 sg13g2_fill_1 FILLER_0_95_804 ();
 sg13g2_fill_2 FILLER_0_95_809 ();
 sg13g2_fill_2 FILLER_0_95_815 ();
 sg13g2_fill_2 FILLER_0_95_821 ();
 sg13g2_fill_4 FILLER_0_95_828 ();
 sg13g2_fill_8 FILLER_0_95_836 ();
 sg13g2_fill_8 FILLER_0_95_844 ();
 sg13g2_fill_8 FILLER_0_95_852 ();
 sg13g2_fill_8 FILLER_0_95_860 ();
 sg13g2_fill_8 FILLER_0_95_868 ();
 sg13g2_fill_8 FILLER_0_95_876 ();
 sg13g2_fill_1 FILLER_0_95_884 ();
 sg13g2_fill_8 FILLER_0_95_890 ();
 sg13g2_fill_8 FILLER_0_95_898 ();
 sg13g2_fill_2 FILLER_0_95_910 ();
 sg13g2_fill_1 FILLER_0_95_912 ();
 sg13g2_fill_8 FILLER_0_95_918 ();
 sg13g2_fill_2 FILLER_0_95_926 ();
 sg13g2_fill_1 FILLER_0_95_928 ();
 sg13g2_fill_8 FILLER_0_95_939 ();
 sg13g2_fill_4 FILLER_0_95_947 ();
 sg13g2_fill_2 FILLER_0_95_951 ();
 sg13g2_fill_1 FILLER_0_95_953 ();
 sg13g2_fill_2 FILLER_0_95_960 ();
 sg13g2_fill_2 FILLER_0_95_968 ();
 sg13g2_fill_2 FILLER_0_95_975 ();
 sg13g2_fill_1 FILLER_0_95_977 ();
 sg13g2_fill_2 FILLER_0_95_983 ();
 sg13g2_fill_1 FILLER_0_95_985 ();
 sg13g2_fill_2 FILLER_0_95_991 ();
 sg13g2_fill_1 FILLER_0_95_993 ();
 sg13g2_fill_2 FILLER_0_95_998 ();
 sg13g2_fill_2 FILLER_0_95_1006 ();
 sg13g2_fill_1 FILLER_0_95_1008 ();
 sg13g2_fill_2 FILLER_0_95_1015 ();
 sg13g2_fill_8 FILLER_0_95_1021 ();
 sg13g2_fill_8 FILLER_0_95_1029 ();
 sg13g2_fill_8 FILLER_0_95_1037 ();
 sg13g2_fill_8 FILLER_0_95_1045 ();
 sg13g2_fill_8 FILLER_0_95_1053 ();
 sg13g2_fill_2 FILLER_0_95_1061 ();
 sg13g2_fill_8 FILLER_0_95_1068 ();
 sg13g2_fill_1 FILLER_0_95_1076 ();
 sg13g2_fill_2 FILLER_0_95_1082 ();
 sg13g2_fill_4 FILLER_0_95_1089 ();
 sg13g2_fill_8 FILLER_0_95_1098 ();
 sg13g2_fill_1 FILLER_0_95_1106 ();
 sg13g2_fill_2 FILLER_0_95_1115 ();
 sg13g2_fill_2 FILLER_0_95_1124 ();
 sg13g2_fill_2 FILLER_0_95_1131 ();
 sg13g2_fill_4 FILLER_0_95_1139 ();
 sg13g2_fill_4 FILLER_0_95_1147 ();
 sg13g2_fill_2 FILLER_0_95_1151 ();
 sg13g2_fill_1 FILLER_0_95_1153 ();
 sg13g2_fill_2 FILLER_0_95_1160 ();
 sg13g2_fill_2 FILLER_0_95_1167 ();
 sg13g2_fill_2 FILLER_0_95_1172 ();
 sg13g2_fill_2 FILLER_0_95_1182 ();
 sg13g2_fill_2 FILLER_0_95_1187 ();
 sg13g2_fill_8 FILLER_0_95_1193 ();
 sg13g2_fill_8 FILLER_0_95_1201 ();
 sg13g2_fill_8 FILLER_0_95_1209 ();
 sg13g2_fill_8 FILLER_0_95_1217 ();
 sg13g2_fill_2 FILLER_0_95_1225 ();
 sg13g2_fill_1 FILLER_0_95_1227 ();
 sg13g2_fill_2 FILLER_0_95_1232 ();
 sg13g2_fill_2 FILLER_0_95_1238 ();
 sg13g2_fill_4 FILLER_0_95_1245 ();
 sg13g2_fill_2 FILLER_0_95_1249 ();
 sg13g2_fill_2 FILLER_0_95_1259 ();
 sg13g2_fill_2 FILLER_0_95_1271 ();
 sg13g2_fill_2 FILLER_0_95_1277 ();
 sg13g2_fill_2 FILLER_0_95_1287 ();
 sg13g2_fill_4 FILLER_0_95_1293 ();
 sg13g2_fill_8 FILLER_0_96_0 ();
 sg13g2_fill_8 FILLER_0_96_8 ();
 sg13g2_fill_8 FILLER_0_96_16 ();
 sg13g2_fill_8 FILLER_0_96_24 ();
 sg13g2_fill_8 FILLER_0_96_32 ();
 sg13g2_fill_8 FILLER_0_96_40 ();
 sg13g2_fill_8 FILLER_0_96_48 ();
 sg13g2_fill_8 FILLER_0_96_56 ();
 sg13g2_fill_8 FILLER_0_96_64 ();
 sg13g2_fill_8 FILLER_0_96_72 ();
 sg13g2_fill_8 FILLER_0_96_80 ();
 sg13g2_fill_8 FILLER_0_96_88 ();
 sg13g2_fill_8 FILLER_0_96_96 ();
 sg13g2_fill_8 FILLER_0_96_104 ();
 sg13g2_fill_8 FILLER_0_96_112 ();
 sg13g2_fill_8 FILLER_0_96_120 ();
 sg13g2_fill_8 FILLER_0_96_128 ();
 sg13g2_fill_8 FILLER_0_96_136 ();
 sg13g2_fill_8 FILLER_0_96_144 ();
 sg13g2_fill_8 FILLER_0_96_152 ();
 sg13g2_fill_8 FILLER_0_96_160 ();
 sg13g2_fill_8 FILLER_0_96_168 ();
 sg13g2_fill_8 FILLER_0_96_176 ();
 sg13g2_fill_8 FILLER_0_96_184 ();
 sg13g2_fill_8 FILLER_0_96_192 ();
 sg13g2_fill_8 FILLER_0_96_200 ();
 sg13g2_fill_8 FILLER_0_96_208 ();
 sg13g2_fill_8 FILLER_0_96_216 ();
 sg13g2_fill_4 FILLER_0_96_224 ();
 sg13g2_fill_2 FILLER_0_96_228 ();
 sg13g2_fill_1 FILLER_0_96_230 ();
 sg13g2_fill_2 FILLER_0_96_257 ();
 sg13g2_fill_2 FILLER_0_96_264 ();
 sg13g2_fill_4 FILLER_0_96_270 ();
 sg13g2_fill_2 FILLER_0_96_274 ();
 sg13g2_fill_1 FILLER_0_96_276 ();
 sg13g2_fill_2 FILLER_0_96_282 ();
 sg13g2_fill_2 FILLER_0_96_290 ();
 sg13g2_fill_2 FILLER_0_96_296 ();
 sg13g2_fill_1 FILLER_0_96_298 ();
 sg13g2_fill_8 FILLER_0_96_304 ();
 sg13g2_fill_8 FILLER_0_96_312 ();
 sg13g2_fill_4 FILLER_0_96_320 ();
 sg13g2_fill_2 FILLER_0_96_324 ();
 sg13g2_fill_2 FILLER_0_96_331 ();
 sg13g2_fill_2 FILLER_0_96_337 ();
 sg13g2_fill_1 FILLER_0_96_339 ();
 sg13g2_fill_2 FILLER_0_96_345 ();
 sg13g2_fill_1 FILLER_0_96_347 ();
 sg13g2_fill_4 FILLER_0_96_358 ();
 sg13g2_fill_1 FILLER_0_96_362 ();
 sg13g2_fill_4 FILLER_0_96_389 ();
 sg13g2_fill_4 FILLER_0_96_398 ();
 sg13g2_fill_1 FILLER_0_96_402 ();
 sg13g2_fill_8 FILLER_0_96_409 ();
 sg13g2_fill_8 FILLER_0_96_417 ();
 sg13g2_fill_2 FILLER_0_96_425 ();
 sg13g2_fill_2 FILLER_0_96_432 ();
 sg13g2_fill_8 FILLER_0_96_442 ();
 sg13g2_fill_8 FILLER_0_96_450 ();
 sg13g2_fill_2 FILLER_0_96_458 ();
 sg13g2_fill_2 FILLER_0_96_465 ();
 sg13g2_fill_8 FILLER_0_96_471 ();
 sg13g2_fill_4 FILLER_0_96_479 ();
 sg13g2_fill_1 FILLER_0_96_483 ();
 sg13g2_fill_2 FILLER_0_96_489 ();
 sg13g2_fill_4 FILLER_0_96_496 ();
 sg13g2_fill_2 FILLER_0_96_505 ();
 sg13g2_fill_2 FILLER_0_96_513 ();
 sg13g2_fill_4 FILLER_0_96_519 ();
 sg13g2_fill_2 FILLER_0_96_523 ();
 sg13g2_fill_1 FILLER_0_96_525 ();
 sg13g2_fill_8 FILLER_0_96_552 ();
 sg13g2_fill_2 FILLER_0_96_560 ();
 sg13g2_fill_8 FILLER_0_96_583 ();
 sg13g2_fill_1 FILLER_0_96_591 ();
 sg13g2_fill_4 FILLER_0_96_597 ();
 sg13g2_fill_2 FILLER_0_96_601 ();
 sg13g2_fill_8 FILLER_0_96_609 ();
 sg13g2_fill_8 FILLER_0_96_617 ();
 sg13g2_fill_4 FILLER_0_96_625 ();
 sg13g2_fill_2 FILLER_0_96_629 ();
 sg13g2_fill_8 FILLER_0_96_657 ();
 sg13g2_fill_4 FILLER_0_96_665 ();
 sg13g2_fill_2 FILLER_0_96_669 ();
 sg13g2_fill_1 FILLER_0_96_671 ();
 sg13g2_fill_4 FILLER_0_96_682 ();
 sg13g2_fill_1 FILLER_0_96_686 ();
 sg13g2_fill_2 FILLER_0_96_713 ();
 sg13g2_fill_8 FILLER_0_96_723 ();
 sg13g2_fill_2 FILLER_0_96_736 ();
 sg13g2_fill_2 FILLER_0_96_743 ();
 sg13g2_fill_1 FILLER_0_96_745 ();
 sg13g2_fill_8 FILLER_0_96_750 ();
 sg13g2_fill_8 FILLER_0_96_758 ();
 sg13g2_fill_8 FILLER_0_96_766 ();
 sg13g2_fill_8 FILLER_0_96_774 ();
 sg13g2_fill_8 FILLER_0_96_782 ();
 sg13g2_fill_4 FILLER_0_96_790 ();
 sg13g2_fill_1 FILLER_0_96_794 ();
 sg13g2_fill_8 FILLER_0_96_800 ();
 sg13g2_fill_2 FILLER_0_96_808 ();
 sg13g2_fill_2 FILLER_0_96_815 ();
 sg13g2_fill_1 FILLER_0_96_817 ();
 sg13g2_fill_8 FILLER_0_96_824 ();
 sg13g2_fill_8 FILLER_0_96_832 ();
 sg13g2_fill_8 FILLER_0_96_840 ();
 sg13g2_fill_8 FILLER_0_96_848 ();
 sg13g2_fill_8 FILLER_0_96_856 ();
 sg13g2_fill_8 FILLER_0_96_864 ();
 sg13g2_fill_8 FILLER_0_96_872 ();
 sg13g2_fill_2 FILLER_0_96_880 ();
 sg13g2_fill_1 FILLER_0_96_882 ();
 sg13g2_fill_8 FILLER_0_96_887 ();
 sg13g2_fill_8 FILLER_0_96_895 ();
 sg13g2_fill_8 FILLER_0_96_903 ();
 sg13g2_fill_2 FILLER_0_96_911 ();
 sg13g2_fill_1 FILLER_0_96_913 ();
 sg13g2_fill_2 FILLER_0_96_919 ();
 sg13g2_fill_8 FILLER_0_96_928 ();
 sg13g2_fill_8 FILLER_0_96_936 ();
 sg13g2_fill_4 FILLER_0_96_944 ();
 sg13g2_fill_2 FILLER_0_96_948 ();
 sg13g2_fill_4 FILLER_0_96_955 ();
 sg13g2_fill_2 FILLER_0_96_959 ();
 sg13g2_fill_2 FILLER_0_96_966 ();
 sg13g2_fill_8 FILLER_0_96_973 ();
 sg13g2_fill_2 FILLER_0_96_981 ();
 sg13g2_fill_2 FILLER_0_96_989 ();
 sg13g2_fill_1 FILLER_0_96_991 ();
 sg13g2_fill_4 FILLER_0_96_1002 ();
 sg13g2_fill_2 FILLER_0_96_1006 ();
 sg13g2_fill_1 FILLER_0_96_1008 ();
 sg13g2_fill_8 FILLER_0_96_1015 ();
 sg13g2_fill_8 FILLER_0_96_1023 ();
 sg13g2_fill_1 FILLER_0_96_1031 ();
 sg13g2_fill_8 FILLER_0_96_1037 ();
 sg13g2_fill_8 FILLER_0_96_1045 ();
 sg13g2_fill_8 FILLER_0_96_1053 ();
 sg13g2_fill_2 FILLER_0_96_1065 ();
 sg13g2_fill_4 FILLER_0_96_1072 ();
 sg13g2_fill_2 FILLER_0_96_1076 ();
 sg13g2_fill_1 FILLER_0_96_1078 ();
 sg13g2_fill_4 FILLER_0_96_1085 ();
 sg13g2_fill_1 FILLER_0_96_1089 ();
 sg13g2_fill_2 FILLER_0_96_1096 ();
 sg13g2_fill_1 FILLER_0_96_1098 ();
 sg13g2_fill_2 FILLER_0_96_1109 ();
 sg13g2_fill_1 FILLER_0_96_1111 ();
 sg13g2_fill_8 FILLER_0_96_1116 ();
 sg13g2_fill_4 FILLER_0_96_1124 ();
 sg13g2_fill_8 FILLER_0_96_1136 ();
 sg13g2_fill_4 FILLER_0_96_1144 ();
 sg13g2_fill_4 FILLER_0_96_1153 ();
 sg13g2_fill_2 FILLER_0_96_1161 ();
 sg13g2_fill_2 FILLER_0_96_1167 ();
 sg13g2_fill_2 FILLER_0_96_1176 ();
 sg13g2_fill_1 FILLER_0_96_1178 ();
 sg13g2_fill_2 FILLER_0_96_1187 ();
 sg13g2_fill_8 FILLER_0_96_1199 ();
 sg13g2_fill_8 FILLER_0_96_1207 ();
 sg13g2_fill_8 FILLER_0_96_1215 ();
 sg13g2_fill_2 FILLER_0_96_1223 ();
 sg13g2_fill_1 FILLER_0_96_1225 ();
 sg13g2_fill_2 FILLER_0_96_1231 ();
 sg13g2_fill_2 FILLER_0_96_1237 ();
 sg13g2_fill_2 FILLER_0_96_1244 ();
 sg13g2_fill_1 FILLER_0_96_1246 ();
 sg13g2_fill_8 FILLER_0_96_1252 ();
 sg13g2_fill_2 FILLER_0_96_1264 ();
 sg13g2_fill_4 FILLER_0_96_1276 ();
 sg13g2_fill_2 FILLER_0_96_1284 ();
 sg13g2_fill_4 FILLER_0_96_1290 ();
 sg13g2_fill_2 FILLER_0_96_1294 ();
 sg13g2_fill_1 FILLER_0_96_1296 ();
 sg13g2_fill_8 FILLER_0_97_0 ();
 sg13g2_fill_8 FILLER_0_97_8 ();
 sg13g2_fill_8 FILLER_0_97_16 ();
 sg13g2_fill_8 FILLER_0_97_24 ();
 sg13g2_fill_8 FILLER_0_97_32 ();
 sg13g2_fill_8 FILLER_0_97_40 ();
 sg13g2_fill_8 FILLER_0_97_48 ();
 sg13g2_fill_8 FILLER_0_97_56 ();
 sg13g2_fill_8 FILLER_0_97_64 ();
 sg13g2_fill_8 FILLER_0_97_72 ();
 sg13g2_fill_8 FILLER_0_97_80 ();
 sg13g2_fill_8 FILLER_0_97_88 ();
 sg13g2_fill_8 FILLER_0_97_96 ();
 sg13g2_fill_8 FILLER_0_97_104 ();
 sg13g2_fill_8 FILLER_0_97_112 ();
 sg13g2_fill_8 FILLER_0_97_120 ();
 sg13g2_fill_8 FILLER_0_97_128 ();
 sg13g2_fill_8 FILLER_0_97_136 ();
 sg13g2_fill_8 FILLER_0_97_144 ();
 sg13g2_fill_8 FILLER_0_97_152 ();
 sg13g2_fill_8 FILLER_0_97_160 ();
 sg13g2_fill_8 FILLER_0_97_168 ();
 sg13g2_fill_8 FILLER_0_97_176 ();
 sg13g2_fill_8 FILLER_0_97_184 ();
 sg13g2_fill_8 FILLER_0_97_192 ();
 sg13g2_fill_8 FILLER_0_97_200 ();
 sg13g2_fill_8 FILLER_0_97_208 ();
 sg13g2_fill_2 FILLER_0_97_242 ();
 sg13g2_fill_4 FILLER_0_97_249 ();
 sg13g2_fill_2 FILLER_0_97_253 ();
 sg13g2_fill_1 FILLER_0_97_255 ();
 sg13g2_fill_2 FILLER_0_97_261 ();
 sg13g2_fill_8 FILLER_0_97_289 ();
 sg13g2_fill_8 FILLER_0_97_297 ();
 sg13g2_fill_4 FILLER_0_97_305 ();
 sg13g2_fill_1 FILLER_0_97_309 ();
 sg13g2_fill_8 FILLER_0_97_318 ();
 sg13g2_fill_2 FILLER_0_97_326 ();
 sg13g2_fill_8 FILLER_0_97_354 ();
 sg13g2_fill_1 FILLER_0_97_362 ();
 sg13g2_fill_8 FILLER_0_97_368 ();
 sg13g2_fill_1 FILLER_0_97_376 ();
 sg13g2_fill_8 FILLER_0_97_382 ();
 sg13g2_fill_8 FILLER_0_97_390 ();
 sg13g2_fill_8 FILLER_0_97_398 ();
 sg13g2_fill_1 FILLER_0_97_406 ();
 sg13g2_fill_8 FILLER_0_97_417 ();
 sg13g2_fill_4 FILLER_0_97_425 ();
 sg13g2_fill_4 FILLER_0_97_434 ();
 sg13g2_fill_1 FILLER_0_97_438 ();
 sg13g2_fill_8 FILLER_0_97_444 ();
 sg13g2_fill_8 FILLER_0_97_452 ();
 sg13g2_fill_2 FILLER_0_97_460 ();
 sg13g2_fill_2 FILLER_0_97_467 ();
 sg13g2_fill_4 FILLER_0_97_474 ();
 sg13g2_fill_1 FILLER_0_97_478 ();
 sg13g2_fill_8 FILLER_0_97_484 ();
 sg13g2_fill_1 FILLER_0_97_492 ();
 sg13g2_fill_8 FILLER_0_97_497 ();
 sg13g2_fill_2 FILLER_0_97_505 ();
 sg13g2_fill_1 FILLER_0_97_507 ();
 sg13g2_fill_2 FILLER_0_97_529 ();
 sg13g2_fill_2 FILLER_0_97_535 ();
 sg13g2_fill_8 FILLER_0_97_542 ();
 sg13g2_fill_1 FILLER_0_97_550 ();
 sg13g2_fill_8 FILLER_0_97_556 ();
 sg13g2_fill_8 FILLER_0_97_564 ();
 sg13g2_fill_4 FILLER_0_97_572 ();
 sg13g2_fill_2 FILLER_0_97_576 ();
 sg13g2_fill_1 FILLER_0_97_578 ();
 sg13g2_fill_2 FILLER_0_97_583 ();
 sg13g2_fill_8 FILLER_0_97_611 ();
 sg13g2_fill_4 FILLER_0_97_619 ();
 sg13g2_fill_1 FILLER_0_97_623 ();
 sg13g2_fill_8 FILLER_0_97_634 ();
 sg13g2_fill_8 FILLER_0_97_642 ();
 sg13g2_fill_8 FILLER_0_97_650 ();
 sg13g2_fill_2 FILLER_0_97_658 ();
 sg13g2_fill_2 FILLER_0_97_681 ();
 sg13g2_fill_2 FILLER_0_97_688 ();
 sg13g2_fill_4 FILLER_0_97_693 ();
 sg13g2_fill_1 FILLER_0_97_697 ();
 sg13g2_fill_8 FILLER_0_97_706 ();
 sg13g2_fill_8 FILLER_0_97_714 ();
 sg13g2_fill_8 FILLER_0_97_722 ();
 sg13g2_fill_2 FILLER_0_97_735 ();
 sg13g2_fill_8 FILLER_0_97_743 ();
 sg13g2_fill_1 FILLER_0_97_751 ();
 sg13g2_fill_8 FILLER_0_97_757 ();
 sg13g2_fill_8 FILLER_0_97_765 ();
 sg13g2_fill_8 FILLER_0_97_773 ();
 sg13g2_fill_8 FILLER_0_97_781 ();
 sg13g2_fill_8 FILLER_0_97_789 ();
 sg13g2_fill_8 FILLER_0_97_801 ();
 sg13g2_fill_4 FILLER_0_97_809 ();
 sg13g2_fill_2 FILLER_0_97_813 ();
 sg13g2_fill_1 FILLER_0_97_815 ();
 sg13g2_fill_8 FILLER_0_97_821 ();
 sg13g2_fill_4 FILLER_0_97_829 ();
 sg13g2_fill_2 FILLER_0_97_833 ();
 sg13g2_fill_8 FILLER_0_97_839 ();
 sg13g2_fill_1 FILLER_0_97_847 ();
 sg13g2_fill_4 FILLER_0_97_853 ();
 sg13g2_fill_2 FILLER_0_97_857 ();
 sg13g2_fill_4 FILLER_0_97_863 ();
 sg13g2_fill_8 FILLER_0_97_871 ();
 sg13g2_fill_8 FILLER_0_97_879 ();
 sg13g2_fill_4 FILLER_0_97_887 ();
 sg13g2_fill_2 FILLER_0_97_891 ();
 sg13g2_fill_1 FILLER_0_97_893 ();
 sg13g2_fill_2 FILLER_0_97_904 ();
 sg13g2_fill_2 FILLER_0_97_911 ();
 sg13g2_fill_2 FILLER_0_97_918 ();
 sg13g2_fill_1 FILLER_0_97_920 ();
 sg13g2_fill_2 FILLER_0_97_926 ();
 sg13g2_fill_8 FILLER_0_97_933 ();
 sg13g2_fill_4 FILLER_0_97_941 ();
 sg13g2_fill_2 FILLER_0_97_945 ();
 sg13g2_fill_1 FILLER_0_97_947 ();
 sg13g2_fill_8 FILLER_0_97_952 ();
 sg13g2_fill_8 FILLER_0_97_960 ();
 sg13g2_fill_8 FILLER_0_97_968 ();
 sg13g2_fill_4 FILLER_0_97_976 ();
 sg13g2_fill_2 FILLER_0_97_985 ();
 sg13g2_fill_4 FILLER_0_97_992 ();
 sg13g2_fill_1 FILLER_0_97_996 ();
 sg13g2_fill_8 FILLER_0_97_1001 ();
 sg13g2_fill_8 FILLER_0_97_1009 ();
 sg13g2_fill_8 FILLER_0_97_1017 ();
 sg13g2_fill_1 FILLER_0_97_1025 ();
 sg13g2_fill_2 FILLER_0_97_1034 ();
 sg13g2_fill_8 FILLER_0_97_1041 ();
 sg13g2_fill_4 FILLER_0_97_1049 ();
 sg13g2_fill_8 FILLER_0_97_1058 ();
 sg13g2_fill_8 FILLER_0_97_1066 ();
 sg13g2_fill_2 FILLER_0_97_1081 ();
 sg13g2_fill_4 FILLER_0_97_1087 ();
 sg13g2_fill_2 FILLER_0_97_1091 ();
 sg13g2_fill_1 FILLER_0_97_1093 ();
 sg13g2_fill_8 FILLER_0_97_1100 ();
 sg13g2_fill_8 FILLER_0_97_1108 ();
 sg13g2_fill_2 FILLER_0_97_1116 ();
 sg13g2_fill_8 FILLER_0_97_1125 ();
 sg13g2_fill_4 FILLER_0_97_1133 ();
 sg13g2_fill_1 FILLER_0_97_1137 ();
 sg13g2_fill_8 FILLER_0_97_1142 ();
 sg13g2_fill_4 FILLER_0_97_1150 ();
 sg13g2_fill_1 FILLER_0_97_1154 ();
 sg13g2_fill_2 FILLER_0_97_1163 ();
 sg13g2_fill_2 FILLER_0_97_1170 ();
 sg13g2_fill_2 FILLER_0_97_1180 ();
 sg13g2_fill_4 FILLER_0_97_1186 ();
 sg13g2_fill_2 FILLER_0_97_1190 ();
 sg13g2_fill_1 FILLER_0_97_1192 ();
 sg13g2_fill_8 FILLER_0_97_1199 ();
 sg13g2_fill_4 FILLER_0_97_1207 ();
 sg13g2_fill_1 FILLER_0_97_1211 ();
 sg13g2_fill_2 FILLER_0_97_1217 ();
 sg13g2_fill_2 FILLER_0_97_1226 ();
 sg13g2_fill_2 FILLER_0_97_1236 ();
 sg13g2_fill_2 FILLER_0_97_1243 ();
 sg13g2_fill_2 FILLER_0_97_1248 ();
 sg13g2_fill_2 FILLER_0_97_1254 ();
 sg13g2_fill_2 FILLER_0_97_1282 ();
 sg13g2_fill_8 FILLER_0_97_1288 ();
 sg13g2_fill_1 FILLER_0_97_1296 ();
 sg13g2_fill_8 FILLER_0_98_0 ();
 sg13g2_fill_8 FILLER_0_98_8 ();
 sg13g2_fill_8 FILLER_0_98_16 ();
 sg13g2_fill_8 FILLER_0_98_24 ();
 sg13g2_fill_8 FILLER_0_98_32 ();
 sg13g2_fill_8 FILLER_0_98_40 ();
 sg13g2_fill_8 FILLER_0_98_48 ();
 sg13g2_fill_8 FILLER_0_98_56 ();
 sg13g2_fill_8 FILLER_0_98_64 ();
 sg13g2_fill_8 FILLER_0_98_72 ();
 sg13g2_fill_8 FILLER_0_98_80 ();
 sg13g2_fill_8 FILLER_0_98_88 ();
 sg13g2_fill_8 FILLER_0_98_96 ();
 sg13g2_fill_8 FILLER_0_98_104 ();
 sg13g2_fill_8 FILLER_0_98_112 ();
 sg13g2_fill_8 FILLER_0_98_120 ();
 sg13g2_fill_8 FILLER_0_98_128 ();
 sg13g2_fill_8 FILLER_0_98_136 ();
 sg13g2_fill_8 FILLER_0_98_144 ();
 sg13g2_fill_8 FILLER_0_98_152 ();
 sg13g2_fill_8 FILLER_0_98_160 ();
 sg13g2_fill_8 FILLER_0_98_168 ();
 sg13g2_fill_8 FILLER_0_98_176 ();
 sg13g2_fill_8 FILLER_0_98_184 ();
 sg13g2_fill_8 FILLER_0_98_192 ();
 sg13g2_fill_8 FILLER_0_98_200 ();
 sg13g2_fill_8 FILLER_0_98_208 ();
 sg13g2_fill_8 FILLER_0_98_216 ();
 sg13g2_fill_8 FILLER_0_98_224 ();
 sg13g2_fill_2 FILLER_0_98_232 ();
 sg13g2_fill_1 FILLER_0_98_234 ();
 sg13g2_fill_2 FILLER_0_98_239 ();
 sg13g2_fill_4 FILLER_0_98_246 ();
 sg13g2_fill_2 FILLER_0_98_250 ();
 sg13g2_fill_2 FILLER_0_98_278 ();
 sg13g2_fill_4 FILLER_0_98_301 ();
 sg13g2_fill_2 FILLER_0_98_305 ();
 sg13g2_fill_2 FILLER_0_98_333 ();
 sg13g2_fill_8 FILLER_0_98_356 ();
 sg13g2_fill_8 FILLER_0_98_364 ();
 sg13g2_fill_4 FILLER_0_98_372 ();
 sg13g2_fill_2 FILLER_0_98_380 ();
 sg13g2_fill_8 FILLER_0_98_408 ();
 sg13g2_fill_4 FILLER_0_98_416 ();
 sg13g2_fill_1 FILLER_0_98_420 ();
 sg13g2_fill_2 FILLER_0_98_426 ();
 sg13g2_fill_2 FILLER_0_98_434 ();
 sg13g2_fill_2 FILLER_0_98_442 ();
 sg13g2_fill_8 FILLER_0_98_448 ();
 sg13g2_fill_8 FILLER_0_98_456 ();
 sg13g2_fill_8 FILLER_0_98_464 ();
 sg13g2_fill_1 FILLER_0_98_472 ();
 sg13g2_fill_8 FILLER_0_98_499 ();
 sg13g2_fill_4 FILLER_0_98_507 ();
 sg13g2_fill_2 FILLER_0_98_511 ();
 sg13g2_fill_1 FILLER_0_98_513 ();
 sg13g2_fill_8 FILLER_0_98_518 ();
 sg13g2_fill_8 FILLER_0_98_526 ();
 sg13g2_fill_2 FILLER_0_98_534 ();
 sg13g2_fill_1 FILLER_0_98_536 ();
 sg13g2_fill_4 FILLER_0_98_542 ();
 sg13g2_fill_2 FILLER_0_98_546 ();
 sg13g2_fill_1 FILLER_0_98_548 ();
 sg13g2_fill_2 FILLER_0_98_553 ();
 sg13g2_fill_1 FILLER_0_98_555 ();
 sg13g2_fill_8 FILLER_0_98_562 ();
 sg13g2_fill_8 FILLER_0_98_570 ();
 sg13g2_fill_2 FILLER_0_98_578 ();
 sg13g2_fill_1 FILLER_0_98_580 ();
 sg13g2_fill_8 FILLER_0_98_586 ();
 sg13g2_fill_2 FILLER_0_98_594 ();
 sg13g2_fill_2 FILLER_0_98_602 ();
 sg13g2_fill_8 FILLER_0_98_608 ();
 sg13g2_fill_8 FILLER_0_98_616 ();
 sg13g2_fill_8 FILLER_0_98_624 ();
 sg13g2_fill_2 FILLER_0_98_642 ();
 sg13g2_fill_8 FILLER_0_98_670 ();
 sg13g2_fill_1 FILLER_0_98_678 ();
 sg13g2_fill_2 FILLER_0_98_684 ();
 sg13g2_fill_2 FILLER_0_98_691 ();
 sg13g2_fill_8 FILLER_0_98_699 ();
 sg13g2_fill_2 FILLER_0_98_707 ();
 sg13g2_fill_8 FILLER_0_98_715 ();
 sg13g2_fill_8 FILLER_0_98_723 ();
 sg13g2_fill_8 FILLER_0_98_731 ();
 sg13g2_fill_4 FILLER_0_98_739 ();
 sg13g2_fill_2 FILLER_0_98_743 ();
 sg13g2_fill_1 FILLER_0_98_745 ();
 sg13g2_fill_8 FILLER_0_98_756 ();
 sg13g2_fill_8 FILLER_0_98_764 ();
 sg13g2_fill_8 FILLER_0_98_777 ();
 sg13g2_fill_4 FILLER_0_98_785 ();
 sg13g2_fill_1 FILLER_0_98_789 ();
 sg13g2_fill_4 FILLER_0_98_794 ();
 sg13g2_fill_1 FILLER_0_98_798 ();
 sg13g2_fill_2 FILLER_0_98_804 ();
 sg13g2_fill_8 FILLER_0_98_813 ();
 sg13g2_fill_8 FILLER_0_98_821 ();
 sg13g2_fill_8 FILLER_0_98_829 ();
 sg13g2_fill_8 FILLER_0_98_837 ();
 sg13g2_fill_2 FILLER_0_98_849 ();
 sg13g2_fill_2 FILLER_0_98_855 ();
 sg13g2_fill_4 FILLER_0_98_863 ();
 sg13g2_fill_1 FILLER_0_98_867 ();
 sg13g2_fill_2 FILLER_0_98_873 ();
 sg13g2_fill_8 FILLER_0_98_880 ();
 sg13g2_fill_8 FILLER_0_98_888 ();
 sg13g2_fill_8 FILLER_0_98_896 ();
 sg13g2_fill_2 FILLER_0_98_904 ();
 sg13g2_fill_2 FILLER_0_98_916 ();
 sg13g2_fill_4 FILLER_0_98_924 ();
 sg13g2_fill_2 FILLER_0_98_928 ();
 sg13g2_fill_1 FILLER_0_98_930 ();
 sg13g2_fill_4 FILLER_0_98_936 ();
 sg13g2_fill_2 FILLER_0_98_940 ();
 sg13g2_fill_2 FILLER_0_98_948 ();
 sg13g2_fill_2 FILLER_0_98_960 ();
 sg13g2_fill_2 FILLER_0_98_968 ();
 sg13g2_fill_8 FILLER_0_98_978 ();
 sg13g2_fill_8 FILLER_0_98_986 ();
 sg13g2_fill_2 FILLER_0_98_994 ();
 sg13g2_fill_8 FILLER_0_98_1001 ();
 sg13g2_fill_8 FILLER_0_98_1009 ();
 sg13g2_fill_2 FILLER_0_98_1017 ();
 sg13g2_fill_8 FILLER_0_98_1023 ();
 sg13g2_fill_8 FILLER_0_98_1031 ();
 sg13g2_fill_8 FILLER_0_98_1039 ();
 sg13g2_fill_4 FILLER_0_98_1047 ();
 sg13g2_fill_2 FILLER_0_98_1051 ();
 sg13g2_fill_1 FILLER_0_98_1053 ();
 sg13g2_fill_2 FILLER_0_98_1061 ();
 sg13g2_fill_4 FILLER_0_98_1069 ();
 sg13g2_fill_2 FILLER_0_98_1073 ();
 sg13g2_fill_1 FILLER_0_98_1075 ();
 sg13g2_fill_8 FILLER_0_98_1084 ();
 sg13g2_fill_8 FILLER_0_98_1100 ();
 sg13g2_fill_4 FILLER_0_98_1108 ();
 sg13g2_fill_2 FILLER_0_98_1112 ();
 sg13g2_fill_1 FILLER_0_98_1114 ();
 sg13g2_fill_2 FILLER_0_98_1121 ();
 sg13g2_fill_4 FILLER_0_98_1131 ();
 sg13g2_fill_1 FILLER_0_98_1135 ();
 sg13g2_fill_4 FILLER_0_98_1140 ();
 sg13g2_fill_1 FILLER_0_98_1144 ();
 sg13g2_fill_4 FILLER_0_98_1150 ();
 sg13g2_fill_2 FILLER_0_98_1160 ();
 sg13g2_fill_2 FILLER_0_98_1167 ();
 sg13g2_fill_2 FILLER_0_98_1177 ();
 sg13g2_fill_4 FILLER_0_98_1184 ();
 sg13g2_fill_2 FILLER_0_98_1188 ();
 sg13g2_fill_1 FILLER_0_98_1190 ();
 sg13g2_fill_8 FILLER_0_98_1195 ();
 sg13g2_fill_8 FILLER_0_98_1203 ();
 sg13g2_fill_8 FILLER_0_98_1211 ();
 sg13g2_fill_8 FILLER_0_98_1219 ();
 sg13g2_fill_4 FILLER_0_98_1227 ();
 sg13g2_fill_1 FILLER_0_98_1231 ();
 sg13g2_fill_8 FILLER_0_98_1237 ();
 sg13g2_fill_8 FILLER_0_98_1245 ();
 sg13g2_fill_2 FILLER_0_98_1253 ();
 sg13g2_fill_2 FILLER_0_98_1265 ();
 sg13g2_fill_2 FILLER_0_98_1271 ();
 sg13g2_fill_8 FILLER_0_98_1277 ();
 sg13g2_fill_2 FILLER_0_98_1285 ();
 sg13g2_fill_4 FILLER_0_98_1291 ();
 sg13g2_fill_2 FILLER_0_98_1295 ();
 sg13g2_fill_8 FILLER_0_99_0 ();
 sg13g2_fill_8 FILLER_0_99_8 ();
 sg13g2_fill_8 FILLER_0_99_16 ();
 sg13g2_fill_8 FILLER_0_99_24 ();
 sg13g2_fill_8 FILLER_0_99_32 ();
 sg13g2_fill_8 FILLER_0_99_40 ();
 sg13g2_fill_8 FILLER_0_99_48 ();
 sg13g2_fill_8 FILLER_0_99_56 ();
 sg13g2_fill_8 FILLER_0_99_64 ();
 sg13g2_fill_8 FILLER_0_99_72 ();
 sg13g2_fill_8 FILLER_0_99_80 ();
 sg13g2_fill_8 FILLER_0_99_88 ();
 sg13g2_fill_8 FILLER_0_99_96 ();
 sg13g2_fill_8 FILLER_0_99_104 ();
 sg13g2_fill_8 FILLER_0_99_112 ();
 sg13g2_fill_8 FILLER_0_99_120 ();
 sg13g2_fill_8 FILLER_0_99_128 ();
 sg13g2_fill_8 FILLER_0_99_136 ();
 sg13g2_fill_8 FILLER_0_99_144 ();
 sg13g2_fill_8 FILLER_0_99_152 ();
 sg13g2_fill_8 FILLER_0_99_160 ();
 sg13g2_fill_8 FILLER_0_99_168 ();
 sg13g2_fill_8 FILLER_0_99_176 ();
 sg13g2_fill_8 FILLER_0_99_184 ();
 sg13g2_fill_8 FILLER_0_99_192 ();
 sg13g2_fill_8 FILLER_0_99_200 ();
 sg13g2_fill_8 FILLER_0_99_208 ();
 sg13g2_fill_8 FILLER_0_99_216 ();
 sg13g2_fill_8 FILLER_0_99_224 ();
 sg13g2_fill_8 FILLER_0_99_232 ();
 sg13g2_fill_8 FILLER_0_99_240 ();
 sg13g2_fill_8 FILLER_0_99_248 ();
 sg13g2_fill_8 FILLER_0_99_256 ();
 sg13g2_fill_8 FILLER_0_99_264 ();
 sg13g2_fill_4 FILLER_0_99_272 ();
 sg13g2_fill_1 FILLER_0_99_276 ();
 sg13g2_fill_8 FILLER_0_99_283 ();
 sg13g2_fill_8 FILLER_0_99_291 ();
 sg13g2_fill_8 FILLER_0_99_299 ();
 sg13g2_fill_4 FILLER_0_99_307 ();
 sg13g2_fill_8 FILLER_0_99_337 ();
 sg13g2_fill_8 FILLER_0_99_345 ();
 sg13g2_fill_8 FILLER_0_99_353 ();
 sg13g2_fill_8 FILLER_0_99_361 ();
 sg13g2_fill_8 FILLER_0_99_369 ();
 sg13g2_fill_8 FILLER_0_99_377 ();
 sg13g2_fill_8 FILLER_0_99_385 ();
 sg13g2_fill_8 FILLER_0_99_393 ();
 sg13g2_fill_8 FILLER_0_99_401 ();
 sg13g2_fill_8 FILLER_0_99_409 ();
 sg13g2_fill_4 FILLER_0_99_417 ();
 sg13g2_fill_1 FILLER_0_99_421 ();
 sg13g2_fill_2 FILLER_0_99_443 ();
 sg13g2_fill_8 FILLER_0_99_471 ();
 sg13g2_fill_8 FILLER_0_99_479 ();
 sg13g2_fill_2 FILLER_0_99_487 ();
 sg13g2_fill_4 FILLER_0_99_494 ();
 sg13g2_fill_1 FILLER_0_99_498 ();
 sg13g2_fill_8 FILLER_0_99_503 ();
 sg13g2_fill_2 FILLER_0_99_511 ();
 sg13g2_fill_2 FILLER_0_99_518 ();
 sg13g2_fill_8 FILLER_0_99_525 ();
 sg13g2_fill_2 FILLER_0_99_538 ();
 sg13g2_fill_8 FILLER_0_99_566 ();
 sg13g2_fill_8 FILLER_0_99_574 ();
 sg13g2_fill_8 FILLER_0_99_582 ();
 sg13g2_fill_1 FILLER_0_99_590 ();
 sg13g2_fill_8 FILLER_0_99_599 ();
 sg13g2_fill_4 FILLER_0_99_607 ();
 sg13g2_fill_2 FILLER_0_99_611 ();
 sg13g2_fill_8 FILLER_0_99_618 ();
 sg13g2_fill_4 FILLER_0_99_626 ();
 sg13g2_fill_2 FILLER_0_99_635 ();
 sg13g2_fill_8 FILLER_0_99_642 ();
 sg13g2_fill_2 FILLER_0_99_650 ();
 sg13g2_fill_2 FILLER_0_99_673 ();
 sg13g2_fill_8 FILLER_0_99_679 ();
 sg13g2_fill_2 FILLER_0_99_687 ();
 sg13g2_fill_4 FILLER_0_99_695 ();
 sg13g2_fill_8 FILLER_0_99_703 ();
 sg13g2_fill_8 FILLER_0_99_711 ();
 sg13g2_fill_4 FILLER_0_99_719 ();
 sg13g2_fill_2 FILLER_0_99_733 ();
 sg13g2_fill_8 FILLER_0_99_761 ();
 sg13g2_fill_1 FILLER_0_99_769 ();
 sg13g2_fill_2 FILLER_0_99_777 ();
 sg13g2_fill_4 FILLER_0_99_805 ();
 sg13g2_fill_2 FILLER_0_99_817 ();
 sg13g2_fill_8 FILLER_0_99_823 ();
 sg13g2_fill_1 FILLER_0_99_831 ();
 sg13g2_fill_2 FILLER_0_99_836 ();
 sg13g2_fill_4 FILLER_0_99_843 ();
 sg13g2_fill_2 FILLER_0_99_847 ();
 sg13g2_fill_1 FILLER_0_99_849 ();
 sg13g2_fill_2 FILLER_0_99_856 ();
 sg13g2_fill_2 FILLER_0_99_865 ();
 sg13g2_fill_8 FILLER_0_99_871 ();
 sg13g2_fill_8 FILLER_0_99_879 ();
 sg13g2_fill_8 FILLER_0_99_887 ();
 sg13g2_fill_8 FILLER_0_99_895 ();
 sg13g2_fill_8 FILLER_0_99_903 ();
 sg13g2_fill_8 FILLER_0_99_911 ();
 sg13g2_fill_8 FILLER_0_99_919 ();
 sg13g2_fill_1 FILLER_0_99_927 ();
 sg13g2_fill_8 FILLER_0_99_932 ();
 sg13g2_fill_8 FILLER_0_99_940 ();
 sg13g2_fill_2 FILLER_0_99_958 ();
 sg13g2_fill_2 FILLER_0_99_966 ();
 sg13g2_fill_2 FILLER_0_99_974 ();
 sg13g2_fill_1 FILLER_0_99_976 ();
 sg13g2_fill_2 FILLER_0_99_987 ();
 sg13g2_fill_8 FILLER_0_99_993 ();
 sg13g2_fill_8 FILLER_0_99_1001 ();
 sg13g2_fill_8 FILLER_0_99_1009 ();
 sg13g2_fill_8 FILLER_0_99_1017 ();
 sg13g2_fill_8 FILLER_0_99_1033 ();
 sg13g2_fill_8 FILLER_0_99_1041 ();
 sg13g2_fill_2 FILLER_0_99_1049 ();
 sg13g2_fill_1 FILLER_0_99_1051 ();
 sg13g2_fill_2 FILLER_0_99_1056 ();
 sg13g2_fill_8 FILLER_0_99_1063 ();
 sg13g2_fill_8 FILLER_0_99_1071 ();
 sg13g2_fill_8 FILLER_0_99_1079 ();
 sg13g2_fill_8 FILLER_0_99_1092 ();
 sg13g2_fill_4 FILLER_0_99_1100 ();
 sg13g2_fill_2 FILLER_0_99_1104 ();
 sg13g2_fill_1 FILLER_0_99_1106 ();
 sg13g2_fill_4 FILLER_0_99_1114 ();
 sg13g2_fill_2 FILLER_0_99_1118 ();
 sg13g2_fill_8 FILLER_0_99_1125 ();
 sg13g2_fill_8 FILLER_0_99_1133 ();
 sg13g2_fill_8 FILLER_0_99_1141 ();
 sg13g2_fill_8 FILLER_0_99_1149 ();
 sg13g2_fill_1 FILLER_0_99_1157 ();
 sg13g2_fill_2 FILLER_0_99_1164 ();
 sg13g2_fill_2 FILLER_0_99_1171 ();
 sg13g2_fill_1 FILLER_0_99_1173 ();
 sg13g2_fill_8 FILLER_0_99_1182 ();
 sg13g2_fill_2 FILLER_0_99_1190 ();
 sg13g2_fill_8 FILLER_0_99_1197 ();
 sg13g2_fill_8 FILLER_0_99_1205 ();
 sg13g2_fill_8 FILLER_0_99_1213 ();
 sg13g2_fill_8 FILLER_0_99_1221 ();
 sg13g2_fill_4 FILLER_0_99_1229 ();
 sg13g2_fill_2 FILLER_0_99_1233 ();
 sg13g2_fill_8 FILLER_0_99_1239 ();
 sg13g2_fill_2 FILLER_0_99_1247 ();
 sg13g2_fill_1 FILLER_0_99_1249 ();
 sg13g2_fill_8 FILLER_0_99_1254 ();
 sg13g2_fill_2 FILLER_0_99_1262 ();
 sg13g2_fill_8 FILLER_0_99_1268 ();
 sg13g2_fill_4 FILLER_0_99_1276 ();
 sg13g2_fill_8 FILLER_0_99_1284 ();
 sg13g2_fill_1 FILLER_0_99_1296 ();
 sg13g2_fill_8 FILLER_0_100_0 ();
 sg13g2_fill_8 FILLER_0_100_8 ();
 sg13g2_fill_8 FILLER_0_100_16 ();
 sg13g2_fill_8 FILLER_0_100_24 ();
 sg13g2_fill_8 FILLER_0_100_32 ();
 sg13g2_fill_8 FILLER_0_100_40 ();
 sg13g2_fill_8 FILLER_0_100_48 ();
 sg13g2_fill_8 FILLER_0_100_56 ();
 sg13g2_fill_8 FILLER_0_100_64 ();
 sg13g2_fill_8 FILLER_0_100_72 ();
 sg13g2_fill_8 FILLER_0_100_80 ();
 sg13g2_fill_8 FILLER_0_100_88 ();
 sg13g2_fill_8 FILLER_0_100_96 ();
 sg13g2_fill_8 FILLER_0_100_104 ();
 sg13g2_fill_8 FILLER_0_100_112 ();
 sg13g2_fill_8 FILLER_0_100_120 ();
 sg13g2_fill_8 FILLER_0_100_128 ();
 sg13g2_fill_8 FILLER_0_100_136 ();
 sg13g2_fill_8 FILLER_0_100_144 ();
 sg13g2_fill_8 FILLER_0_100_152 ();
 sg13g2_fill_8 FILLER_0_100_160 ();
 sg13g2_fill_8 FILLER_0_100_168 ();
 sg13g2_fill_8 FILLER_0_100_176 ();
 sg13g2_fill_8 FILLER_0_100_184 ();
 sg13g2_fill_8 FILLER_0_100_192 ();
 sg13g2_fill_8 FILLER_0_100_200 ();
 sg13g2_fill_8 FILLER_0_100_208 ();
 sg13g2_fill_8 FILLER_0_100_216 ();
 sg13g2_fill_8 FILLER_0_100_224 ();
 sg13g2_fill_8 FILLER_0_100_232 ();
 sg13g2_fill_8 FILLER_0_100_240 ();
 sg13g2_fill_8 FILLER_0_100_248 ();
 sg13g2_fill_8 FILLER_0_100_256 ();
 sg13g2_fill_8 FILLER_0_100_264 ();
 sg13g2_fill_8 FILLER_0_100_272 ();
 sg13g2_fill_4 FILLER_0_100_280 ();
 sg13g2_fill_1 FILLER_0_100_284 ();
 sg13g2_fill_4 FILLER_0_100_291 ();
 sg13g2_fill_2 FILLER_0_100_295 ();
 sg13g2_fill_2 FILLER_0_100_302 ();
 sg13g2_fill_4 FILLER_0_100_309 ();
 sg13g2_fill_8 FILLER_0_100_317 ();
 sg13g2_fill_4 FILLER_0_100_325 ();
 sg13g2_fill_2 FILLER_0_100_339 ();
 sg13g2_fill_2 FILLER_0_100_345 ();
 sg13g2_fill_4 FILLER_0_100_352 ();
 sg13g2_fill_1 FILLER_0_100_356 ();
 sg13g2_fill_8 FILLER_0_100_361 ();
 sg13g2_fill_8 FILLER_0_100_390 ();
 sg13g2_fill_2 FILLER_0_100_398 ();
 sg13g2_fill_2 FILLER_0_100_410 ();
 sg13g2_fill_2 FILLER_0_100_417 ();
 sg13g2_fill_1 FILLER_0_100_419 ();
 sg13g2_fill_4 FILLER_0_100_424 ();
 sg13g2_fill_8 FILLER_0_100_432 ();
 sg13g2_fill_4 FILLER_0_100_440 ();
 sg13g2_fill_1 FILLER_0_100_444 ();
 sg13g2_fill_8 FILLER_0_100_450 ();
 sg13g2_fill_4 FILLER_0_100_458 ();
 sg13g2_fill_8 FILLER_0_100_466 ();
 sg13g2_fill_8 FILLER_0_100_474 ();
 sg13g2_fill_8 FILLER_0_100_482 ();
 sg13g2_fill_8 FILLER_0_100_490 ();
 sg13g2_fill_4 FILLER_0_100_498 ();
 sg13g2_fill_2 FILLER_0_100_502 ();
 sg13g2_fill_2 FILLER_0_100_509 ();
 sg13g2_fill_8 FILLER_0_100_537 ();
 sg13g2_fill_8 FILLER_0_100_545 ();
 sg13g2_fill_1 FILLER_0_100_553 ();
 sg13g2_fill_2 FILLER_0_100_559 ();
 sg13g2_fill_2 FILLER_0_100_587 ();
 sg13g2_fill_1 FILLER_0_100_589 ();
 sg13g2_fill_8 FILLER_0_100_596 ();
 sg13g2_fill_8 FILLER_0_100_604 ();
 sg13g2_fill_8 FILLER_0_100_612 ();
 sg13g2_fill_2 FILLER_0_100_620 ();
 sg13g2_fill_1 FILLER_0_100_622 ();
 sg13g2_fill_4 FILLER_0_100_633 ();
 sg13g2_fill_2 FILLER_0_100_642 ();
 sg13g2_fill_1 FILLER_0_100_644 ();
 sg13g2_fill_2 FILLER_0_100_649 ();
 sg13g2_fill_8 FILLER_0_100_656 ();
 sg13g2_fill_2 FILLER_0_100_674 ();
 sg13g2_fill_8 FILLER_0_100_702 ();
 sg13g2_fill_1 FILLER_0_100_710 ();
 sg13g2_fill_4 FILLER_0_100_715 ();
 sg13g2_fill_2 FILLER_0_100_724 ();
 sg13g2_fill_2 FILLER_0_100_752 ();
 sg13g2_fill_4 FILLER_0_100_759 ();
 sg13g2_fill_8 FILLER_0_100_767 ();
 sg13g2_fill_2 FILLER_0_100_780 ();
 sg13g2_fill_2 FILLER_0_100_792 ();
 sg13g2_fill_8 FILLER_0_100_798 ();
 sg13g2_fill_8 FILLER_0_100_806 ();
 sg13g2_fill_1 FILLER_0_100_814 ();
 sg13g2_fill_4 FILLER_0_100_819 ();
 sg13g2_fill_1 FILLER_0_100_823 ();
 sg13g2_fill_4 FILLER_0_100_830 ();
 sg13g2_fill_1 FILLER_0_100_834 ();
 sg13g2_fill_8 FILLER_0_100_840 ();
 sg13g2_fill_8 FILLER_0_100_848 ();
 sg13g2_fill_4 FILLER_0_100_856 ();
 sg13g2_fill_8 FILLER_0_100_865 ();
 sg13g2_fill_1 FILLER_0_100_873 ();
 sg13g2_fill_8 FILLER_0_100_879 ();
 sg13g2_fill_8 FILLER_0_100_887 ();
 sg13g2_fill_8 FILLER_0_100_895 ();
 sg13g2_fill_4 FILLER_0_100_903 ();
 sg13g2_fill_8 FILLER_0_100_912 ();
 sg13g2_fill_8 FILLER_0_100_920 ();
 sg13g2_fill_8 FILLER_0_100_928 ();
 sg13g2_fill_1 FILLER_0_100_936 ();
 sg13g2_fill_8 FILLER_0_100_941 ();
 sg13g2_fill_8 FILLER_0_100_949 ();
 sg13g2_fill_4 FILLER_0_100_957 ();
 sg13g2_fill_8 FILLER_0_100_967 ();
 sg13g2_fill_2 FILLER_0_100_975 ();
 sg13g2_fill_1 FILLER_0_100_977 ();
 sg13g2_fill_2 FILLER_0_100_982 ();
 sg13g2_fill_4 FILLER_0_100_989 ();
 sg13g2_fill_1 FILLER_0_100_993 ();
 sg13g2_fill_2 FILLER_0_100_998 ();
 sg13g2_fill_2 FILLER_0_100_1005 ();
 sg13g2_fill_1 FILLER_0_100_1007 ();
 sg13g2_fill_2 FILLER_0_100_1013 ();
 sg13g2_fill_8 FILLER_0_100_1023 ();
 sg13g2_fill_8 FILLER_0_100_1031 ();
 sg13g2_fill_8 FILLER_0_100_1039 ();
 sg13g2_fill_8 FILLER_0_100_1047 ();
 sg13g2_fill_2 FILLER_0_100_1060 ();
 sg13g2_fill_8 FILLER_0_100_1068 ();
 sg13g2_fill_8 FILLER_0_100_1076 ();
 sg13g2_fill_8 FILLER_0_100_1094 ();
 sg13g2_fill_4 FILLER_0_100_1102 ();
 sg13g2_fill_2 FILLER_0_100_1106 ();
 sg13g2_fill_2 FILLER_0_100_1115 ();
 sg13g2_fill_2 FILLER_0_100_1125 ();
 sg13g2_fill_8 FILLER_0_100_1132 ();
 sg13g2_fill_8 FILLER_0_100_1140 ();
 sg13g2_fill_8 FILLER_0_100_1148 ();
 sg13g2_fill_1 FILLER_0_100_1156 ();
 sg13g2_fill_2 FILLER_0_100_1162 ();
 sg13g2_fill_8 FILLER_0_100_1171 ();
 sg13g2_fill_2 FILLER_0_100_1184 ();
 sg13g2_fill_1 FILLER_0_100_1186 ();
 sg13g2_fill_2 FILLER_0_100_1191 ();
 sg13g2_fill_8 FILLER_0_100_1198 ();
 sg13g2_fill_8 FILLER_0_100_1206 ();
 sg13g2_fill_8 FILLER_0_100_1214 ();
 sg13g2_fill_2 FILLER_0_100_1227 ();
 sg13g2_fill_2 FILLER_0_100_1234 ();
 sg13g2_fill_8 FILLER_0_100_1241 ();
 sg13g2_fill_8 FILLER_0_100_1249 ();
 sg13g2_fill_4 FILLER_0_100_1257 ();
 sg13g2_fill_2 FILLER_0_100_1261 ();
 sg13g2_fill_1 FILLER_0_100_1263 ();
 sg13g2_fill_4 FILLER_0_100_1268 ();
 sg13g2_fill_1 FILLER_0_100_1272 ();
 sg13g2_fill_2 FILLER_0_100_1277 ();
 sg13g2_fill_8 FILLER_0_100_1284 ();
 sg13g2_fill_4 FILLER_0_100_1292 ();
 sg13g2_fill_1 FILLER_0_100_1296 ();
 sg13g2_fill_8 FILLER_0_101_0 ();
 sg13g2_fill_8 FILLER_0_101_8 ();
 sg13g2_fill_8 FILLER_0_101_16 ();
 sg13g2_fill_8 FILLER_0_101_24 ();
 sg13g2_fill_8 FILLER_0_101_32 ();
 sg13g2_fill_8 FILLER_0_101_40 ();
 sg13g2_fill_8 FILLER_0_101_48 ();
 sg13g2_fill_8 FILLER_0_101_56 ();
 sg13g2_fill_8 FILLER_0_101_64 ();
 sg13g2_fill_8 FILLER_0_101_72 ();
 sg13g2_fill_8 FILLER_0_101_80 ();
 sg13g2_fill_8 FILLER_0_101_88 ();
 sg13g2_fill_8 FILLER_0_101_96 ();
 sg13g2_fill_8 FILLER_0_101_104 ();
 sg13g2_fill_8 FILLER_0_101_112 ();
 sg13g2_fill_8 FILLER_0_101_120 ();
 sg13g2_fill_8 FILLER_0_101_128 ();
 sg13g2_fill_8 FILLER_0_101_136 ();
 sg13g2_fill_8 FILLER_0_101_144 ();
 sg13g2_fill_8 FILLER_0_101_152 ();
 sg13g2_fill_8 FILLER_0_101_160 ();
 sg13g2_fill_8 FILLER_0_101_168 ();
 sg13g2_fill_8 FILLER_0_101_176 ();
 sg13g2_fill_8 FILLER_0_101_184 ();
 sg13g2_fill_8 FILLER_0_101_192 ();
 sg13g2_fill_8 FILLER_0_101_200 ();
 sg13g2_fill_8 FILLER_0_101_208 ();
 sg13g2_fill_2 FILLER_0_101_216 ();
 sg13g2_fill_1 FILLER_0_101_218 ();
 sg13g2_fill_2 FILLER_0_101_245 ();
 sg13g2_fill_2 FILLER_0_101_251 ();
 sg13g2_fill_4 FILLER_0_101_279 ();
 sg13g2_fill_2 FILLER_0_101_293 ();
 sg13g2_fill_8 FILLER_0_101_300 ();
 sg13g2_fill_8 FILLER_0_101_308 ();
 sg13g2_fill_1 FILLER_0_101_316 ();
 sg13g2_fill_2 FILLER_0_101_322 ();
 sg13g2_fill_8 FILLER_0_101_328 ();
 sg13g2_fill_8 FILLER_0_101_336 ();
 sg13g2_fill_1 FILLER_0_101_344 ();
 sg13g2_fill_2 FILLER_0_101_350 ();
 sg13g2_fill_4 FILLER_0_101_378 ();
 sg13g2_fill_2 FILLER_0_101_382 ();
 sg13g2_fill_2 FILLER_0_101_389 ();
 sg13g2_fill_8 FILLER_0_101_395 ();
 sg13g2_fill_4 FILLER_0_101_403 ();
 sg13g2_fill_8 FILLER_0_101_433 ();
 sg13g2_fill_4 FILLER_0_101_441 ();
 sg13g2_fill_1 FILLER_0_101_445 ();
 sg13g2_fill_8 FILLER_0_101_450 ();
 sg13g2_fill_8 FILLER_0_101_458 ();
 sg13g2_fill_8 FILLER_0_101_466 ();
 sg13g2_fill_8 FILLER_0_101_474 ();
 sg13g2_fill_8 FILLER_0_101_482 ();
 sg13g2_fill_1 FILLER_0_101_490 ();
 sg13g2_fill_8 FILLER_0_101_517 ();
 sg13g2_fill_8 FILLER_0_101_525 ();
 sg13g2_fill_8 FILLER_0_101_533 ();
 sg13g2_fill_8 FILLER_0_101_541 ();
 sg13g2_fill_8 FILLER_0_101_549 ();
 sg13g2_fill_8 FILLER_0_101_557 ();
 sg13g2_fill_4 FILLER_0_101_570 ();
 sg13g2_fill_1 FILLER_0_101_574 ();
 sg13g2_fill_8 FILLER_0_101_579 ();
 sg13g2_fill_8 FILLER_0_101_587 ();
 sg13g2_fill_1 FILLER_0_101_595 ();
 sg13g2_fill_8 FILLER_0_101_602 ();
 sg13g2_fill_2 FILLER_0_101_610 ();
 sg13g2_fill_1 FILLER_0_101_612 ();
 sg13g2_fill_8 FILLER_0_101_618 ();
 sg13g2_fill_4 FILLER_0_101_626 ();
 sg13g2_fill_8 FILLER_0_101_656 ();
 sg13g2_fill_4 FILLER_0_101_664 ();
 sg13g2_fill_8 FILLER_0_101_672 ();
 sg13g2_fill_8 FILLER_0_101_680 ();
 sg13g2_fill_2 FILLER_0_101_688 ();
 sg13g2_fill_1 FILLER_0_101_690 ();
 sg13g2_fill_8 FILLER_0_101_696 ();
 sg13g2_fill_4 FILLER_0_101_704 ();
 sg13g2_fill_1 FILLER_0_101_708 ();
 sg13g2_fill_4 FILLER_0_101_714 ();
 sg13g2_fill_2 FILLER_0_101_718 ();
 sg13g2_fill_1 FILLER_0_101_720 ();
 sg13g2_fill_8 FILLER_0_101_731 ();
 sg13g2_fill_4 FILLER_0_101_739 ();
 sg13g2_fill_4 FILLER_0_101_753 ();
 sg13g2_fill_2 FILLER_0_101_757 ();
 sg13g2_fill_8 FILLER_0_101_769 ();
 sg13g2_fill_8 FILLER_0_101_777 ();
 sg13g2_fill_8 FILLER_0_101_785 ();
 sg13g2_fill_2 FILLER_0_101_793 ();
 sg13g2_fill_1 FILLER_0_101_795 ();
 sg13g2_fill_8 FILLER_0_101_801 ();
 sg13g2_fill_2 FILLER_0_101_809 ();
 sg13g2_fill_2 FILLER_0_101_821 ();
 sg13g2_fill_4 FILLER_0_101_827 ();
 sg13g2_fill_2 FILLER_0_101_831 ();
 sg13g2_fill_2 FILLER_0_101_843 ();
 sg13g2_fill_4 FILLER_0_101_850 ();
 sg13g2_fill_2 FILLER_0_101_854 ();
 sg13g2_fill_4 FILLER_0_101_861 ();
 sg13g2_fill_8 FILLER_0_101_870 ();
 sg13g2_fill_4 FILLER_0_101_878 ();
 sg13g2_fill_1 FILLER_0_101_882 ();
 sg13g2_fill_2 FILLER_0_101_904 ();
 sg13g2_fill_8 FILLER_0_101_927 ();
 sg13g2_fill_4 FILLER_0_101_935 ();
 sg13g2_fill_2 FILLER_0_101_944 ();
 sg13g2_fill_4 FILLER_0_101_950 ();
 sg13g2_fill_2 FILLER_0_101_954 ();
 sg13g2_fill_2 FILLER_0_101_963 ();
 sg13g2_fill_2 FILLER_0_101_969 ();
 sg13g2_fill_4 FILLER_0_101_976 ();
 sg13g2_fill_1 FILLER_0_101_980 ();
 sg13g2_fill_8 FILLER_0_101_986 ();
 sg13g2_fill_4 FILLER_0_101_994 ();
 sg13g2_fill_2 FILLER_0_101_998 ();
 sg13g2_fill_8 FILLER_0_101_1005 ();
 sg13g2_fill_2 FILLER_0_101_1013 ();
 sg13g2_fill_2 FILLER_0_101_1019 ();
 sg13g2_fill_1 FILLER_0_101_1021 ();
 sg13g2_fill_8 FILLER_0_101_1027 ();
 sg13g2_fill_1 FILLER_0_101_1035 ();
 sg13g2_fill_8 FILLER_0_101_1041 ();
 sg13g2_fill_4 FILLER_0_101_1049 ();
 sg13g2_fill_2 FILLER_0_101_1053 ();
 sg13g2_fill_4 FILLER_0_101_1059 ();
 sg13g2_fill_1 FILLER_0_101_1063 ();
 sg13g2_fill_2 FILLER_0_101_1068 ();
 sg13g2_fill_4 FILLER_0_101_1078 ();
 sg13g2_fill_2 FILLER_0_101_1082 ();
 sg13g2_fill_1 FILLER_0_101_1084 ();
 sg13g2_fill_2 FILLER_0_101_1089 ();
 sg13g2_fill_8 FILLER_0_101_1096 ();
 sg13g2_fill_8 FILLER_0_101_1104 ();
 sg13g2_fill_4 FILLER_0_101_1112 ();
 sg13g2_fill_2 FILLER_0_101_1123 ();
 sg13g2_fill_8 FILLER_0_101_1130 ();
 sg13g2_fill_8 FILLER_0_101_1138 ();
 sg13g2_fill_8 FILLER_0_101_1146 ();
 sg13g2_fill_8 FILLER_0_101_1154 ();
 sg13g2_fill_8 FILLER_0_101_1162 ();
 sg13g2_fill_2 FILLER_0_101_1170 ();
 sg13g2_fill_1 FILLER_0_101_1172 ();
 sg13g2_fill_8 FILLER_0_101_1178 ();
 sg13g2_fill_1 FILLER_0_101_1186 ();
 sg13g2_fill_8 FILLER_0_101_1192 ();
 sg13g2_fill_8 FILLER_0_101_1200 ();
 sg13g2_fill_8 FILLER_0_101_1208 ();
 sg13g2_fill_8 FILLER_0_101_1216 ();
 sg13g2_fill_1 FILLER_0_101_1224 ();
 sg13g2_fill_2 FILLER_0_101_1232 ();
 sg13g2_fill_2 FILLER_0_101_1241 ();
 sg13g2_fill_2 FILLER_0_101_1248 ();
 sg13g2_fill_2 FILLER_0_101_1276 ();
 sg13g2_fill_8 FILLER_0_101_1285 ();
 sg13g2_fill_4 FILLER_0_101_1293 ();
 sg13g2_fill_8 FILLER_0_102_0 ();
 sg13g2_fill_8 FILLER_0_102_8 ();
 sg13g2_fill_8 FILLER_0_102_16 ();
 sg13g2_fill_8 FILLER_0_102_24 ();
 sg13g2_fill_8 FILLER_0_102_32 ();
 sg13g2_fill_8 FILLER_0_102_40 ();
 sg13g2_fill_8 FILLER_0_102_48 ();
 sg13g2_fill_8 FILLER_0_102_56 ();
 sg13g2_fill_8 FILLER_0_102_64 ();
 sg13g2_fill_8 FILLER_0_102_72 ();
 sg13g2_fill_8 FILLER_0_102_80 ();
 sg13g2_fill_8 FILLER_0_102_88 ();
 sg13g2_fill_8 FILLER_0_102_96 ();
 sg13g2_fill_8 FILLER_0_102_104 ();
 sg13g2_fill_8 FILLER_0_102_112 ();
 sg13g2_fill_8 FILLER_0_102_120 ();
 sg13g2_fill_8 FILLER_0_102_128 ();
 sg13g2_fill_8 FILLER_0_102_136 ();
 sg13g2_fill_8 FILLER_0_102_144 ();
 sg13g2_fill_8 FILLER_0_102_152 ();
 sg13g2_fill_8 FILLER_0_102_160 ();
 sg13g2_fill_8 FILLER_0_102_168 ();
 sg13g2_fill_8 FILLER_0_102_176 ();
 sg13g2_fill_8 FILLER_0_102_184 ();
 sg13g2_fill_8 FILLER_0_102_192 ();
 sg13g2_fill_8 FILLER_0_102_200 ();
 sg13g2_fill_8 FILLER_0_102_208 ();
 sg13g2_fill_2 FILLER_0_102_216 ();
 sg13g2_fill_1 FILLER_0_102_218 ();
 sg13g2_fill_4 FILLER_0_102_224 ();
 sg13g2_fill_4 FILLER_0_102_254 ();
 sg13g2_fill_2 FILLER_0_102_258 ();
 sg13g2_fill_4 FILLER_0_102_265 ();
 sg13g2_fill_2 FILLER_0_102_269 ();
 sg13g2_fill_4 FILLER_0_102_292 ();
 sg13g2_fill_1 FILLER_0_102_296 ();
 sg13g2_fill_8 FILLER_0_102_301 ();
 sg13g2_fill_8 FILLER_0_102_309 ();
 sg13g2_fill_8 FILLER_0_102_317 ();
 sg13g2_fill_8 FILLER_0_102_325 ();
 sg13g2_fill_4 FILLER_0_102_333 ();
 sg13g2_fill_1 FILLER_0_102_337 ();
 sg13g2_fill_8 FILLER_0_102_343 ();
 sg13g2_fill_8 FILLER_0_102_351 ();
 sg13g2_fill_4 FILLER_0_102_359 ();
 sg13g2_fill_2 FILLER_0_102_363 ();
 sg13g2_fill_1 FILLER_0_102_365 ();
 sg13g2_fill_8 FILLER_0_102_392 ();
 sg13g2_fill_8 FILLER_0_102_400 ();
 sg13g2_fill_8 FILLER_0_102_408 ();
 sg13g2_fill_2 FILLER_0_102_421 ();
 sg13g2_fill_1 FILLER_0_102_423 ();
 sg13g2_fill_2 FILLER_0_102_429 ();
 sg13g2_fill_4 FILLER_0_102_437 ();
 sg13g2_fill_1 FILLER_0_102_441 ();
 sg13g2_fill_4 FILLER_0_102_454 ();
 sg13g2_fill_2 FILLER_0_102_458 ();
 sg13g2_fill_1 FILLER_0_102_460 ();
 sg13g2_fill_4 FILLER_0_102_466 ();
 sg13g2_fill_2 FILLER_0_102_475 ();
 sg13g2_fill_8 FILLER_0_102_481 ();
 sg13g2_fill_8 FILLER_0_102_489 ();
 sg13g2_fill_8 FILLER_0_102_497 ();
 sg13g2_fill_8 FILLER_0_102_505 ();
 sg13g2_fill_8 FILLER_0_102_513 ();
 sg13g2_fill_8 FILLER_0_102_521 ();
 sg13g2_fill_8 FILLER_0_102_529 ();
 sg13g2_fill_8 FILLER_0_102_537 ();
 sg13g2_fill_8 FILLER_0_102_545 ();
 sg13g2_fill_8 FILLER_0_102_553 ();
 sg13g2_fill_8 FILLER_0_102_561 ();
 sg13g2_fill_8 FILLER_0_102_569 ();
 sg13g2_fill_8 FILLER_0_102_577 ();
 sg13g2_fill_8 FILLER_0_102_585 ();
 sg13g2_fill_2 FILLER_0_102_593 ();
 sg13g2_fill_8 FILLER_0_102_600 ();
 sg13g2_fill_8 FILLER_0_102_608 ();
 sg13g2_fill_8 FILLER_0_102_616 ();
 sg13g2_fill_2 FILLER_0_102_624 ();
 sg13g2_fill_2 FILLER_0_102_636 ();
 sg13g2_fill_8 FILLER_0_102_642 ();
 sg13g2_fill_8 FILLER_0_102_650 ();
 sg13g2_fill_4 FILLER_0_102_658 ();
 sg13g2_fill_1 FILLER_0_102_662 ();
 sg13g2_fill_2 FILLER_0_102_689 ();
 sg13g2_fill_2 FILLER_0_102_712 ();
 sg13g2_fill_8 FILLER_0_102_724 ();
 sg13g2_fill_4 FILLER_0_102_732 ();
 sg13g2_fill_8 FILLER_0_102_746 ();
 sg13g2_fill_8 FILLER_0_102_754 ();
 sg13g2_fill_4 FILLER_0_102_762 ();
 sg13g2_fill_2 FILLER_0_102_766 ();
 sg13g2_fill_1 FILLER_0_102_768 ();
 sg13g2_fill_8 FILLER_0_102_775 ();
 sg13g2_fill_8 FILLER_0_102_783 ();
 sg13g2_fill_2 FILLER_0_102_791 ();
 sg13g2_fill_1 FILLER_0_102_793 ();
 sg13g2_fill_8 FILLER_0_102_799 ();
 sg13g2_fill_4 FILLER_0_102_807 ();
 sg13g2_fill_1 FILLER_0_102_811 ();
 sg13g2_fill_2 FILLER_0_102_822 ();
 sg13g2_fill_2 FILLER_0_102_828 ();
 sg13g2_fill_2 FILLER_0_102_856 ();
 sg13g2_fill_8 FILLER_0_102_862 ();
 sg13g2_fill_8 FILLER_0_102_870 ();
 sg13g2_fill_2 FILLER_0_102_878 ();
 sg13g2_fill_1 FILLER_0_102_880 ();
 sg13g2_fill_2 FILLER_0_102_902 ();
 sg13g2_fill_2 FILLER_0_102_925 ();
 sg13g2_fill_8 FILLER_0_102_932 ();
 sg13g2_fill_2 FILLER_0_102_940 ();
 sg13g2_fill_1 FILLER_0_102_942 ();
 sg13g2_fill_2 FILLER_0_102_948 ();
 sg13g2_fill_2 FILLER_0_102_956 ();
 sg13g2_fill_4 FILLER_0_102_963 ();
 sg13g2_fill_1 FILLER_0_102_967 ();
 sg13g2_fill_2 FILLER_0_102_974 ();
 sg13g2_fill_4 FILLER_0_102_980 ();
 sg13g2_fill_2 FILLER_0_102_984 ();
 sg13g2_fill_8 FILLER_0_102_990 ();
 sg13g2_fill_8 FILLER_0_102_998 ();
 sg13g2_fill_2 FILLER_0_102_1014 ();
 sg13g2_fill_2 FILLER_0_102_1021 ();
 sg13g2_fill_8 FILLER_0_102_1029 ();
 sg13g2_fill_8 FILLER_0_102_1037 ();
 sg13g2_fill_8 FILLER_0_102_1045 ();
 sg13g2_fill_2 FILLER_0_102_1057 ();
 sg13g2_fill_2 FILLER_0_102_1064 ();
 sg13g2_fill_8 FILLER_0_102_1071 ();
 sg13g2_fill_8 FILLER_0_102_1079 ();
 sg13g2_fill_2 FILLER_0_102_1087 ();
 sg13g2_fill_2 FILLER_0_102_1099 ();
 sg13g2_fill_4 FILLER_0_102_1109 ();
 sg13g2_fill_2 FILLER_0_102_1113 ();
 sg13g2_fill_1 FILLER_0_102_1115 ();
 sg13g2_fill_2 FILLER_0_102_1121 ();
 sg13g2_fill_8 FILLER_0_102_1131 ();
 sg13g2_fill_8 FILLER_0_102_1139 ();
 sg13g2_fill_2 FILLER_0_102_1147 ();
 sg13g2_fill_1 FILLER_0_102_1149 ();
 sg13g2_fill_8 FILLER_0_102_1154 ();
 sg13g2_fill_2 FILLER_0_102_1162 ();
 sg13g2_fill_2 FILLER_0_102_1168 ();
 sg13g2_fill_4 FILLER_0_102_1175 ();
 sg13g2_fill_1 FILLER_0_102_1179 ();
 sg13g2_fill_4 FILLER_0_102_1186 ();
 sg13g2_fill_2 FILLER_0_102_1190 ();
 sg13g2_fill_1 FILLER_0_102_1192 ();
 sg13g2_fill_8 FILLER_0_102_1199 ();
 sg13g2_fill_8 FILLER_0_102_1207 ();
 sg13g2_fill_1 FILLER_0_102_1215 ();
 sg13g2_fill_4 FILLER_0_102_1224 ();
 sg13g2_fill_1 FILLER_0_102_1228 ();
 sg13g2_fill_2 FILLER_0_102_1234 ();
 sg13g2_fill_2 FILLER_0_102_1244 ();
 sg13g2_fill_1 FILLER_0_102_1246 ();
 sg13g2_fill_2 FILLER_0_102_1255 ();
 sg13g2_fill_4 FILLER_0_102_1262 ();
 sg13g2_fill_1 FILLER_0_102_1266 ();
 sg13g2_fill_4 FILLER_0_102_1273 ();
 sg13g2_fill_1 FILLER_0_102_1277 ();
 sg13g2_fill_4 FILLER_0_102_1282 ();
 sg13g2_fill_1 FILLER_0_102_1286 ();
 sg13g2_fill_4 FILLER_0_102_1291 ();
 sg13g2_fill_2 FILLER_0_102_1295 ();
 sg13g2_fill_8 FILLER_0_103_0 ();
 sg13g2_fill_8 FILLER_0_103_8 ();
 sg13g2_fill_8 FILLER_0_103_16 ();
 sg13g2_fill_8 FILLER_0_103_24 ();
 sg13g2_fill_8 FILLER_0_103_32 ();
 sg13g2_fill_8 FILLER_0_103_40 ();
 sg13g2_fill_8 FILLER_0_103_48 ();
 sg13g2_fill_8 FILLER_0_103_56 ();
 sg13g2_fill_8 FILLER_0_103_64 ();
 sg13g2_fill_8 FILLER_0_103_72 ();
 sg13g2_fill_8 FILLER_0_103_80 ();
 sg13g2_fill_8 FILLER_0_103_88 ();
 sg13g2_fill_8 FILLER_0_103_96 ();
 sg13g2_fill_8 FILLER_0_103_104 ();
 sg13g2_fill_8 FILLER_0_103_112 ();
 sg13g2_fill_8 FILLER_0_103_120 ();
 sg13g2_fill_8 FILLER_0_103_128 ();
 sg13g2_fill_8 FILLER_0_103_136 ();
 sg13g2_fill_8 FILLER_0_103_144 ();
 sg13g2_fill_8 FILLER_0_103_152 ();
 sg13g2_fill_8 FILLER_0_103_160 ();
 sg13g2_fill_8 FILLER_0_103_168 ();
 sg13g2_fill_8 FILLER_0_103_176 ();
 sg13g2_fill_8 FILLER_0_103_184 ();
 sg13g2_fill_8 FILLER_0_103_192 ();
 sg13g2_fill_8 FILLER_0_103_200 ();
 sg13g2_fill_8 FILLER_0_103_208 ();
 sg13g2_fill_8 FILLER_0_103_216 ();
 sg13g2_fill_2 FILLER_0_103_228 ();
 sg13g2_fill_1 FILLER_0_103_230 ();
 sg13g2_fill_2 FILLER_0_103_236 ();
 sg13g2_fill_1 FILLER_0_103_238 ();
 sg13g2_fill_4 FILLER_0_103_244 ();
 sg13g2_fill_4 FILLER_0_103_254 ();
 sg13g2_fill_4 FILLER_0_103_263 ();
 sg13g2_fill_1 FILLER_0_103_267 ();
 sg13g2_fill_2 FILLER_0_103_294 ();
 sg13g2_fill_8 FILLER_0_103_301 ();
 sg13g2_fill_8 FILLER_0_103_309 ();
 sg13g2_fill_8 FILLER_0_103_317 ();
 sg13g2_fill_8 FILLER_0_103_325 ();
 sg13g2_fill_2 FILLER_0_103_333 ();
 sg13g2_fill_1 FILLER_0_103_335 ();
 sg13g2_fill_2 FILLER_0_103_362 ();
 sg13g2_fill_1 FILLER_0_103_364 ();
 sg13g2_fill_8 FILLER_0_103_386 ();
 sg13g2_fill_8 FILLER_0_103_394 ();
 sg13g2_fill_2 FILLER_0_103_402 ();
 sg13g2_fill_8 FILLER_0_103_409 ();
 sg13g2_fill_8 FILLER_0_103_417 ();
 sg13g2_fill_2 FILLER_0_103_425 ();
 sg13g2_fill_1 FILLER_0_103_427 ();
 sg13g2_fill_2 FILLER_0_103_434 ();
 sg13g2_fill_2 FILLER_0_103_441 ();
 sg13g2_fill_2 FILLER_0_103_449 ();
 sg13g2_fill_4 FILLER_0_103_457 ();
 sg13g2_fill_2 FILLER_0_103_466 ();
 sg13g2_fill_2 FILLER_0_103_494 ();
 sg13g2_fill_4 FILLER_0_103_501 ();
 sg13g2_fill_2 FILLER_0_103_510 ();
 sg13g2_fill_8 FILLER_0_103_516 ();
 sg13g2_fill_8 FILLER_0_103_524 ();
 sg13g2_fill_8 FILLER_0_103_532 ();
 sg13g2_fill_2 FILLER_0_103_540 ();
 sg13g2_fill_4 FILLER_0_103_547 ();
 sg13g2_fill_2 FILLER_0_103_551 ();
 sg13g2_fill_1 FILLER_0_103_553 ();
 sg13g2_fill_4 FILLER_0_103_558 ();
 sg13g2_fill_1 FILLER_0_103_562 ();
 sg13g2_fill_2 FILLER_0_103_567 ();
 sg13g2_fill_2 FILLER_0_103_574 ();
 sg13g2_fill_4 FILLER_0_103_602 ();
 sg13g2_fill_2 FILLER_0_103_606 ();
 sg13g2_fill_8 FILLER_0_103_613 ();
 sg13g2_fill_1 FILLER_0_103_621 ();
 sg13g2_fill_4 FILLER_0_103_648 ();
 sg13g2_fill_2 FILLER_0_103_652 ();
 sg13g2_fill_1 FILLER_0_103_654 ();
 sg13g2_fill_8 FILLER_0_103_665 ();
 sg13g2_fill_4 FILLER_0_103_673 ();
 sg13g2_fill_1 FILLER_0_103_677 ();
 sg13g2_fill_4 FILLER_0_103_683 ();
 sg13g2_fill_2 FILLER_0_103_692 ();
 sg13g2_fill_1 FILLER_0_103_694 ();
 sg13g2_fill_2 FILLER_0_103_701 ();
 sg13g2_fill_1 FILLER_0_103_703 ();
 sg13g2_fill_4 FILLER_0_103_730 ();
 sg13g2_fill_8 FILLER_0_103_760 ();
 sg13g2_fill_4 FILLER_0_103_768 ();
 sg13g2_fill_1 FILLER_0_103_772 ();
 sg13g2_fill_2 FILLER_0_103_779 ();
 sg13g2_fill_2 FILLER_0_103_789 ();
 sg13g2_fill_8 FILLER_0_103_798 ();
 sg13g2_fill_2 FILLER_0_103_806 ();
 sg13g2_fill_1 FILLER_0_103_808 ();
 sg13g2_fill_2 FILLER_0_103_814 ();
 sg13g2_fill_8 FILLER_0_103_842 ();
 sg13g2_fill_4 FILLER_0_103_850 ();
 sg13g2_fill_8 FILLER_0_103_858 ();
 sg13g2_fill_8 FILLER_0_103_866 ();
 sg13g2_fill_8 FILLER_0_103_874 ();
 sg13g2_fill_8 FILLER_0_103_882 ();
 sg13g2_fill_8 FILLER_0_103_890 ();
 sg13g2_fill_1 FILLER_0_103_898 ();
 sg13g2_fill_2 FILLER_0_103_904 ();
 sg13g2_fill_2 FILLER_0_103_927 ();
 sg13g2_fill_8 FILLER_0_103_950 ();
 sg13g2_fill_8 FILLER_0_103_958 ();
 sg13g2_fill_8 FILLER_0_103_966 ();
 sg13g2_fill_4 FILLER_0_103_974 ();
 sg13g2_fill_2 FILLER_0_103_983 ();
 sg13g2_fill_8 FILLER_0_103_990 ();
 sg13g2_fill_8 FILLER_0_103_998 ();
 sg13g2_fill_1 FILLER_0_103_1006 ();
 sg13g2_fill_2 FILLER_0_103_1012 ();
 sg13g2_fill_8 FILLER_0_103_1019 ();
 sg13g2_fill_8 FILLER_0_103_1027 ();
 sg13g2_fill_8 FILLER_0_103_1035 ();
 sg13g2_fill_4 FILLER_0_103_1043 ();
 sg13g2_fill_2 FILLER_0_103_1047 ();
 sg13g2_fill_8 FILLER_0_103_1057 ();
 sg13g2_fill_8 FILLER_0_103_1065 ();
 sg13g2_fill_4 FILLER_0_103_1073 ();
 sg13g2_fill_1 FILLER_0_103_1077 ();
 sg13g2_fill_4 FILLER_0_103_1082 ();
 sg13g2_fill_2 FILLER_0_103_1086 ();
 sg13g2_fill_1 FILLER_0_103_1088 ();
 sg13g2_fill_2 FILLER_0_103_1093 ();
 sg13g2_fill_8 FILLER_0_103_1100 ();
 sg13g2_fill_8 FILLER_0_103_1108 ();
 sg13g2_fill_2 FILLER_0_103_1116 ();
 sg13g2_fill_1 FILLER_0_103_1118 ();
 sg13g2_fill_2 FILLER_0_103_1124 ();
 sg13g2_fill_2 FILLER_0_103_1131 ();
 sg13g2_fill_2 FILLER_0_103_1137 ();
 sg13g2_fill_1 FILLER_0_103_1139 ();
 sg13g2_fill_2 FILLER_0_103_1145 ();
 sg13g2_fill_1 FILLER_0_103_1147 ();
 sg13g2_fill_2 FILLER_0_103_1154 ();
 sg13g2_fill_1 FILLER_0_103_1156 ();
 sg13g2_fill_2 FILLER_0_103_1165 ();
 sg13g2_fill_2 FILLER_0_103_1172 ();
 sg13g2_fill_2 FILLER_0_103_1180 ();
 sg13g2_fill_2 FILLER_0_103_1189 ();
 sg13g2_fill_2 FILLER_0_103_1196 ();
 sg13g2_fill_8 FILLER_0_103_1203 ();
 sg13g2_fill_8 FILLER_0_103_1211 ();
 sg13g2_fill_2 FILLER_0_103_1219 ();
 sg13g2_fill_1 FILLER_0_103_1221 ();
 sg13g2_fill_2 FILLER_0_103_1227 ();
 sg13g2_fill_4 FILLER_0_103_1236 ();
 sg13g2_fill_2 FILLER_0_103_1247 ();
 sg13g2_fill_8 FILLER_0_103_1254 ();
 sg13g2_fill_2 FILLER_0_103_1262 ();
 sg13g2_fill_1 FILLER_0_103_1264 ();
 sg13g2_fill_8 FILLER_0_103_1269 ();
 sg13g2_fill_4 FILLER_0_103_1281 ();
 sg13g2_fill_4 FILLER_0_103_1290 ();
 sg13g2_fill_2 FILLER_0_103_1294 ();
 sg13g2_fill_1 FILLER_0_103_1296 ();
 sg13g2_fill_8 FILLER_0_104_0 ();
 sg13g2_fill_8 FILLER_0_104_8 ();
 sg13g2_fill_8 FILLER_0_104_16 ();
 sg13g2_fill_8 FILLER_0_104_24 ();
 sg13g2_fill_8 FILLER_0_104_32 ();
 sg13g2_fill_8 FILLER_0_104_40 ();
 sg13g2_fill_8 FILLER_0_104_48 ();
 sg13g2_fill_8 FILLER_0_104_56 ();
 sg13g2_fill_8 FILLER_0_104_64 ();
 sg13g2_fill_8 FILLER_0_104_72 ();
 sg13g2_fill_8 FILLER_0_104_80 ();
 sg13g2_fill_8 FILLER_0_104_88 ();
 sg13g2_fill_8 FILLER_0_104_96 ();
 sg13g2_fill_8 FILLER_0_104_104 ();
 sg13g2_fill_8 FILLER_0_104_112 ();
 sg13g2_fill_8 FILLER_0_104_120 ();
 sg13g2_fill_8 FILLER_0_104_128 ();
 sg13g2_fill_8 FILLER_0_104_136 ();
 sg13g2_fill_8 FILLER_0_104_144 ();
 sg13g2_fill_8 FILLER_0_104_152 ();
 sg13g2_fill_8 FILLER_0_104_160 ();
 sg13g2_fill_8 FILLER_0_104_168 ();
 sg13g2_fill_8 FILLER_0_104_176 ();
 sg13g2_fill_8 FILLER_0_104_184 ();
 sg13g2_fill_8 FILLER_0_104_192 ();
 sg13g2_fill_8 FILLER_0_104_200 ();
 sg13g2_fill_8 FILLER_0_104_208 ();
 sg13g2_fill_8 FILLER_0_104_216 ();
 sg13g2_fill_8 FILLER_0_104_224 ();
 sg13g2_fill_8 FILLER_0_104_232 ();
 sg13g2_fill_4 FILLER_0_104_240 ();
 sg13g2_fill_2 FILLER_0_104_244 ();
 sg13g2_fill_8 FILLER_0_104_250 ();
 sg13g2_fill_2 FILLER_0_104_258 ();
 sg13g2_fill_8 FILLER_0_104_264 ();
 sg13g2_fill_8 FILLER_0_104_272 ();
 sg13g2_fill_4 FILLER_0_104_280 ();
 sg13g2_fill_2 FILLER_0_104_284 ();
 sg13g2_fill_1 FILLER_0_104_286 ();
 sg13g2_fill_2 FILLER_0_104_292 ();
 sg13g2_fill_8 FILLER_0_104_320 ();
 sg13g2_fill_8 FILLER_0_104_328 ();
 sg13g2_fill_8 FILLER_0_104_336 ();
 sg13g2_fill_4 FILLER_0_104_344 ();
 sg13g2_fill_2 FILLER_0_104_348 ();
 sg13g2_fill_1 FILLER_0_104_350 ();
 sg13g2_fill_2 FILLER_0_104_355 ();
 sg13g2_fill_8 FILLER_0_104_361 ();
 sg13g2_fill_2 FILLER_0_104_369 ();
 sg13g2_fill_2 FILLER_0_104_381 ();
 sg13g2_fill_8 FILLER_0_104_388 ();
 sg13g2_fill_8 FILLER_0_104_396 ();
 sg13g2_fill_8 FILLER_0_104_404 ();
 sg13g2_fill_8 FILLER_0_104_417 ();
 sg13g2_fill_2 FILLER_0_104_425 ();
 sg13g2_fill_8 FILLER_0_104_432 ();
 sg13g2_fill_4 FILLER_0_104_440 ();
 sg13g2_fill_1 FILLER_0_104_444 ();
 sg13g2_fill_8 FILLER_0_104_453 ();
 sg13g2_fill_4 FILLER_0_104_461 ();
 sg13g2_fill_2 FILLER_0_104_465 ();
 sg13g2_fill_2 FILLER_0_104_472 ();
 sg13g2_fill_8 FILLER_0_104_478 ();
 sg13g2_fill_1 FILLER_0_104_486 ();
 sg13g2_fill_4 FILLER_0_104_492 ();
 sg13g2_fill_2 FILLER_0_104_496 ();
 sg13g2_fill_2 FILLER_0_104_524 ();
 sg13g2_fill_4 FILLER_0_104_531 ();
 sg13g2_fill_2 FILLER_0_104_535 ();
 sg13g2_fill_1 FILLER_0_104_537 ();
 sg13g2_fill_2 FILLER_0_104_564 ();
 sg13g2_fill_8 FILLER_0_104_576 ();
 sg13g2_fill_8 FILLER_0_104_584 ();
 sg13g2_fill_2 FILLER_0_104_592 ();
 sg13g2_fill_8 FILLER_0_104_599 ();
 sg13g2_fill_8 FILLER_0_104_607 ();
 sg13g2_fill_4 FILLER_0_104_615 ();
 sg13g2_fill_2 FILLER_0_104_619 ();
 sg13g2_fill_8 FILLER_0_104_626 ();
 sg13g2_fill_8 FILLER_0_104_634 ();
 sg13g2_fill_4 FILLER_0_104_642 ();
 sg13g2_fill_2 FILLER_0_104_646 ();
 sg13g2_fill_1 FILLER_0_104_648 ();
 sg13g2_fill_2 FILLER_0_104_653 ();
 sg13g2_fill_2 FILLER_0_104_681 ();
 sg13g2_fill_8 FILLER_0_104_688 ();
 sg13g2_fill_1 FILLER_0_104_696 ();
 sg13g2_fill_8 FILLER_0_104_707 ();
 sg13g2_fill_8 FILLER_0_104_715 ();
 sg13g2_fill_2 FILLER_0_104_723 ();
 sg13g2_fill_1 FILLER_0_104_725 ();
 sg13g2_fill_4 FILLER_0_104_752 ();
 sg13g2_fill_2 FILLER_0_104_766 ();
 sg13g2_fill_4 FILLER_0_104_773 ();
 sg13g2_fill_2 FILLER_0_104_777 ();
 sg13g2_fill_4 FILLER_0_104_784 ();
 sg13g2_fill_1 FILLER_0_104_788 ();
 sg13g2_fill_2 FILLER_0_104_794 ();
 sg13g2_fill_2 FILLER_0_104_801 ();
 sg13g2_fill_2 FILLER_0_104_808 ();
 sg13g2_fill_8 FILLER_0_104_814 ();
 sg13g2_fill_4 FILLER_0_104_822 ();
 sg13g2_fill_4 FILLER_0_104_831 ();
 sg13g2_fill_1 FILLER_0_104_835 ();
 sg13g2_fill_4 FILLER_0_104_846 ();
 sg13g2_fill_2 FILLER_0_104_850 ();
 sg13g2_fill_1 FILLER_0_104_852 ();
 sg13g2_fill_2 FILLER_0_104_858 ();
 sg13g2_fill_2 FILLER_0_104_867 ();
 sg13g2_fill_1 FILLER_0_104_869 ();
 sg13g2_fill_2 FILLER_0_104_875 ();
 sg13g2_fill_2 FILLER_0_104_883 ();
 sg13g2_fill_8 FILLER_0_104_889 ();
 sg13g2_fill_1 FILLER_0_104_897 ();
 sg13g2_fill_8 FILLER_0_104_902 ();
 sg13g2_fill_8 FILLER_0_104_910 ();
 sg13g2_fill_8 FILLER_0_104_918 ();
 sg13g2_fill_4 FILLER_0_104_926 ();
 sg13g2_fill_2 FILLER_0_104_930 ();
 sg13g2_fill_2 FILLER_0_104_937 ();
 sg13g2_fill_8 FILLER_0_104_946 ();
 sg13g2_fill_8 FILLER_0_104_954 ();
 sg13g2_fill_4 FILLER_0_104_962 ();
 sg13g2_fill_1 FILLER_0_104_966 ();
 sg13g2_fill_2 FILLER_0_104_972 ();
 sg13g2_fill_1 FILLER_0_104_974 ();
 sg13g2_fill_4 FILLER_0_104_979 ();
 sg13g2_fill_2 FILLER_0_104_989 ();
 sg13g2_fill_1 FILLER_0_104_991 ();
 sg13g2_fill_4 FILLER_0_104_999 ();
 sg13g2_fill_8 FILLER_0_104_1011 ();
 sg13g2_fill_8 FILLER_0_104_1019 ();
 sg13g2_fill_8 FILLER_0_104_1027 ();
 sg13g2_fill_4 FILLER_0_104_1035 ();
 sg13g2_fill_2 FILLER_0_104_1039 ();
 sg13g2_fill_2 FILLER_0_104_1046 ();
 sg13g2_fill_4 FILLER_0_104_1056 ();
 sg13g2_fill_2 FILLER_0_104_1060 ();
 sg13g2_fill_1 FILLER_0_104_1062 ();
 sg13g2_fill_4 FILLER_0_104_1067 ();
 sg13g2_fill_2 FILLER_0_104_1071 ();
 sg13g2_fill_8 FILLER_0_104_1081 ();
 sg13g2_fill_4 FILLER_0_104_1089 ();
 sg13g2_fill_2 FILLER_0_104_1093 ();
 sg13g2_fill_4 FILLER_0_104_1100 ();
 sg13g2_fill_2 FILLER_0_104_1109 ();
 sg13g2_fill_1 FILLER_0_104_1111 ();
 sg13g2_fill_8 FILLER_0_104_1116 ();
 sg13g2_fill_1 FILLER_0_104_1124 ();
 sg13g2_fill_2 FILLER_0_104_1130 ();
 sg13g2_fill_1 FILLER_0_104_1132 ();
 sg13g2_fill_4 FILLER_0_104_1138 ();
 sg13g2_fill_2 FILLER_0_104_1142 ();
 sg13g2_fill_1 FILLER_0_104_1144 ();
 sg13g2_fill_8 FILLER_0_104_1148 ();
 sg13g2_fill_2 FILLER_0_104_1160 ();
 sg13g2_fill_4 FILLER_0_104_1167 ();
 sg13g2_fill_1 FILLER_0_104_1171 ();
 sg13g2_fill_2 FILLER_0_104_1177 ();
 sg13g2_fill_2 FILLER_0_104_1184 ();
 sg13g2_fill_2 FILLER_0_104_1191 ();
 sg13g2_fill_1 FILLER_0_104_1193 ();
 sg13g2_fill_8 FILLER_0_104_1200 ();
 sg13g2_fill_8 FILLER_0_104_1208 ();
 sg13g2_fill_4 FILLER_0_104_1216 ();
 sg13g2_fill_2 FILLER_0_104_1220 ();
 sg13g2_fill_1 FILLER_0_104_1222 ();
 sg13g2_fill_8 FILLER_0_104_1228 ();
 sg13g2_fill_4 FILLER_0_104_1236 ();
 sg13g2_fill_1 FILLER_0_104_1240 ();
 sg13g2_fill_8 FILLER_0_104_1249 ();
 sg13g2_fill_8 FILLER_0_104_1257 ();
 sg13g2_fill_8 FILLER_0_104_1265 ();
 sg13g2_fill_2 FILLER_0_104_1281 ();
 sg13g2_fill_2 FILLER_0_104_1287 ();
 sg13g2_fill_4 FILLER_0_104_1293 ();
 sg13g2_fill_8 FILLER_0_105_0 ();
 sg13g2_fill_8 FILLER_0_105_8 ();
 sg13g2_fill_8 FILLER_0_105_16 ();
 sg13g2_fill_8 FILLER_0_105_24 ();
 sg13g2_fill_8 FILLER_0_105_32 ();
 sg13g2_fill_8 FILLER_0_105_40 ();
 sg13g2_fill_8 FILLER_0_105_48 ();
 sg13g2_fill_8 FILLER_0_105_56 ();
 sg13g2_fill_8 FILLER_0_105_64 ();
 sg13g2_fill_8 FILLER_0_105_72 ();
 sg13g2_fill_8 FILLER_0_105_80 ();
 sg13g2_fill_8 FILLER_0_105_88 ();
 sg13g2_fill_8 FILLER_0_105_96 ();
 sg13g2_fill_8 FILLER_0_105_104 ();
 sg13g2_fill_8 FILLER_0_105_112 ();
 sg13g2_fill_8 FILLER_0_105_120 ();
 sg13g2_fill_8 FILLER_0_105_128 ();
 sg13g2_fill_8 FILLER_0_105_136 ();
 sg13g2_fill_8 FILLER_0_105_144 ();
 sg13g2_fill_8 FILLER_0_105_152 ();
 sg13g2_fill_8 FILLER_0_105_160 ();
 sg13g2_fill_8 FILLER_0_105_168 ();
 sg13g2_fill_8 FILLER_0_105_176 ();
 sg13g2_fill_8 FILLER_0_105_184 ();
 sg13g2_fill_8 FILLER_0_105_192 ();
 sg13g2_fill_8 FILLER_0_105_200 ();
 sg13g2_fill_8 FILLER_0_105_208 ();
 sg13g2_fill_8 FILLER_0_105_216 ();
 sg13g2_fill_8 FILLER_0_105_224 ();
 sg13g2_fill_8 FILLER_0_105_232 ();
 sg13g2_fill_8 FILLER_0_105_240 ();
 sg13g2_fill_8 FILLER_0_105_248 ();
 sg13g2_fill_4 FILLER_0_105_256 ();
 sg13g2_fill_8 FILLER_0_105_265 ();
 sg13g2_fill_8 FILLER_0_105_273 ();
 sg13g2_fill_8 FILLER_0_105_281 ();
 sg13g2_fill_2 FILLER_0_105_289 ();
 sg13g2_fill_1 FILLER_0_105_291 ();
 sg13g2_fill_2 FILLER_0_105_296 ();
 sg13g2_fill_2 FILLER_0_105_303 ();
 sg13g2_fill_2 FILLER_0_105_310 ();
 sg13g2_fill_8 FILLER_0_105_316 ();
 sg13g2_fill_2 FILLER_0_105_324 ();
 sg13g2_fill_1 FILLER_0_105_326 ();
 sg13g2_fill_8 FILLER_0_105_331 ();
 sg13g2_fill_4 FILLER_0_105_339 ();
 sg13g2_fill_2 FILLER_0_105_343 ();
 sg13g2_fill_1 FILLER_0_105_345 ();
 sg13g2_fill_2 FILLER_0_105_351 ();
 sg13g2_fill_8 FILLER_0_105_379 ();
 sg13g2_fill_8 FILLER_0_105_391 ();
 sg13g2_fill_2 FILLER_0_105_399 ();
 sg13g2_fill_1 FILLER_0_105_401 ();
 sg13g2_fill_2 FILLER_0_105_428 ();
 sg13g2_fill_8 FILLER_0_105_435 ();
 sg13g2_fill_4 FILLER_0_105_443 ();
 sg13g2_fill_2 FILLER_0_105_447 ();
 sg13g2_fill_2 FILLER_0_105_454 ();
 sg13g2_fill_8 FILLER_0_105_477 ();
 sg13g2_fill_8 FILLER_0_105_485 ();
 sg13g2_fill_1 FILLER_0_105_493 ();
 sg13g2_fill_8 FILLER_0_105_499 ();
 sg13g2_fill_8 FILLER_0_105_507 ();
 sg13g2_fill_2 FILLER_0_105_515 ();
 sg13g2_fill_2 FILLER_0_105_527 ();
 sg13g2_fill_8 FILLER_0_105_555 ();
 sg13g2_fill_2 FILLER_0_105_563 ();
 sg13g2_fill_1 FILLER_0_105_565 ();
 sg13g2_fill_2 FILLER_0_105_569 ();
 sg13g2_fill_2 FILLER_0_105_575 ();
 sg13g2_fill_2 FILLER_0_105_583 ();
 sg13g2_fill_2 FILLER_0_105_593 ();
 sg13g2_fill_8 FILLER_0_105_600 ();
 sg13g2_fill_4 FILLER_0_105_608 ();
 sg13g2_fill_8 FILLER_0_105_617 ();
 sg13g2_fill_8 FILLER_0_105_625 ();
 sg13g2_fill_8 FILLER_0_105_633 ();
 sg13g2_fill_8 FILLER_0_105_641 ();
 sg13g2_fill_4 FILLER_0_105_649 ();
 sg13g2_fill_1 FILLER_0_105_653 ();
 sg13g2_fill_2 FILLER_0_105_661 ();
 sg13g2_fill_2 FILLER_0_105_668 ();
 sg13g2_fill_8 FILLER_0_105_678 ();
 sg13g2_fill_4 FILLER_0_105_686 ();
 sg13g2_fill_2 FILLER_0_105_690 ();
 sg13g2_fill_1 FILLER_0_105_692 ();
 sg13g2_fill_8 FILLER_0_105_698 ();
 sg13g2_fill_8 FILLER_0_105_706 ();
 sg13g2_fill_8 FILLER_0_105_714 ();
 sg13g2_fill_8 FILLER_0_105_722 ();
 sg13g2_fill_8 FILLER_0_105_730 ();
 sg13g2_fill_2 FILLER_0_105_738 ();
 sg13g2_fill_2 FILLER_0_105_744 ();
 sg13g2_fill_2 FILLER_0_105_750 ();
 sg13g2_fill_8 FILLER_0_105_757 ();
 sg13g2_fill_2 FILLER_0_105_765 ();
 sg13g2_fill_8 FILLER_0_105_793 ();
 sg13g2_fill_8 FILLER_0_105_801 ();
 sg13g2_fill_8 FILLER_0_105_809 ();
 sg13g2_fill_8 FILLER_0_105_817 ();
 sg13g2_fill_8 FILLER_0_105_825 ();
 sg13g2_fill_8 FILLER_0_105_833 ();
 sg13g2_fill_8 FILLER_0_105_841 ();
 sg13g2_fill_8 FILLER_0_105_849 ();
 sg13g2_fill_8 FILLER_0_105_857 ();
 sg13g2_fill_8 FILLER_0_105_865 ();
 sg13g2_fill_8 FILLER_0_105_873 ();
 sg13g2_fill_8 FILLER_0_105_881 ();
 sg13g2_fill_8 FILLER_0_105_889 ();
 sg13g2_fill_8 FILLER_0_105_903 ();
 sg13g2_fill_8 FILLER_0_105_911 ();
 sg13g2_fill_4 FILLER_0_105_919 ();
 sg13g2_fill_2 FILLER_0_105_923 ();
 sg13g2_fill_8 FILLER_0_105_930 ();
 sg13g2_fill_1 FILLER_0_105_938 ();
 sg13g2_fill_2 FILLER_0_105_949 ();
 sg13g2_fill_4 FILLER_0_105_955 ();
 sg13g2_fill_2 FILLER_0_105_959 ();
 sg13g2_fill_1 FILLER_0_105_961 ();
 sg13g2_fill_8 FILLER_0_105_968 ();
 sg13g2_fill_8 FILLER_0_105_976 ();
 sg13g2_fill_2 FILLER_0_105_990 ();
 sg13g2_fill_4 FILLER_0_105_997 ();
 sg13g2_fill_2 FILLER_0_105_1001 ();
 sg13g2_fill_1 FILLER_0_105_1003 ();
 sg13g2_fill_2 FILLER_0_105_1008 ();
 sg13g2_fill_8 FILLER_0_105_1015 ();
 sg13g2_fill_4 FILLER_0_105_1023 ();
 sg13g2_fill_4 FILLER_0_105_1035 ();
 sg13g2_fill_2 FILLER_0_105_1044 ();
 sg13g2_fill_1 FILLER_0_105_1046 ();
 sg13g2_fill_4 FILLER_0_105_1052 ();
 sg13g2_fill_4 FILLER_0_105_1060 ();
 sg13g2_fill_2 FILLER_0_105_1069 ();
 sg13g2_fill_8 FILLER_0_105_1075 ();
 sg13g2_fill_8 FILLER_0_105_1083 ();
 sg13g2_fill_1 FILLER_0_105_1091 ();
 sg13g2_fill_2 FILLER_0_105_1097 ();
 sg13g2_fill_2 FILLER_0_105_1103 ();
 sg13g2_fill_1 FILLER_0_105_1105 ();
 sg13g2_fill_2 FILLER_0_105_1114 ();
 sg13g2_fill_2 FILLER_0_105_1120 ();
 sg13g2_fill_1 FILLER_0_105_1122 ();
 sg13g2_fill_4 FILLER_0_105_1128 ();
 sg13g2_fill_2 FILLER_0_105_1132 ();
 sg13g2_fill_1 FILLER_0_105_1134 ();
 sg13g2_fill_2 FILLER_0_105_1140 ();
 sg13g2_fill_1 FILLER_0_105_1142 ();
 sg13g2_fill_4 FILLER_0_105_1149 ();
 sg13g2_fill_4 FILLER_0_105_1157 ();
 sg13g2_fill_1 FILLER_0_105_1161 ();
 sg13g2_fill_8 FILLER_0_105_1166 ();
 sg13g2_fill_8 FILLER_0_105_1174 ();
 sg13g2_fill_4 FILLER_0_105_1185 ();
 sg13g2_fill_2 FILLER_0_105_1189 ();
 sg13g2_fill_4 FILLER_0_105_1195 ();
 sg13g2_fill_2 FILLER_0_105_1199 ();
 sg13g2_fill_8 FILLER_0_105_1206 ();
 sg13g2_fill_2 FILLER_0_105_1218 ();
 sg13g2_fill_8 FILLER_0_105_1225 ();
 sg13g2_fill_8 FILLER_0_105_1233 ();
 sg13g2_fill_4 FILLER_0_105_1246 ();
 sg13g2_fill_4 FILLER_0_105_1254 ();
 sg13g2_fill_1 FILLER_0_105_1258 ();
 sg13g2_fill_4 FILLER_0_105_1266 ();
 sg13g2_fill_2 FILLER_0_105_1270 ();
 sg13g2_fill_1 FILLER_0_105_1272 ();
 sg13g2_fill_2 FILLER_0_105_1278 ();
 sg13g2_fill_2 FILLER_0_105_1284 ();
 sg13g2_fill_2 FILLER_0_105_1290 ();
 sg13g2_fill_1 FILLER_0_105_1296 ();
 sg13g2_fill_8 FILLER_0_106_0 ();
 sg13g2_fill_8 FILLER_0_106_8 ();
 sg13g2_fill_8 FILLER_0_106_16 ();
 sg13g2_fill_8 FILLER_0_106_24 ();
 sg13g2_fill_8 FILLER_0_106_32 ();
 sg13g2_fill_8 FILLER_0_106_40 ();
 sg13g2_fill_8 FILLER_0_106_48 ();
 sg13g2_fill_8 FILLER_0_106_56 ();
 sg13g2_fill_8 FILLER_0_106_64 ();
 sg13g2_fill_8 FILLER_0_106_72 ();
 sg13g2_fill_8 FILLER_0_106_80 ();
 sg13g2_fill_8 FILLER_0_106_88 ();
 sg13g2_fill_8 FILLER_0_106_96 ();
 sg13g2_fill_8 FILLER_0_106_104 ();
 sg13g2_fill_8 FILLER_0_106_112 ();
 sg13g2_fill_8 FILLER_0_106_120 ();
 sg13g2_fill_8 FILLER_0_106_128 ();
 sg13g2_fill_8 FILLER_0_106_136 ();
 sg13g2_fill_8 FILLER_0_106_144 ();
 sg13g2_fill_8 FILLER_0_106_152 ();
 sg13g2_fill_8 FILLER_0_106_160 ();
 sg13g2_fill_8 FILLER_0_106_168 ();
 sg13g2_fill_8 FILLER_0_106_176 ();
 sg13g2_fill_8 FILLER_0_106_184 ();
 sg13g2_fill_8 FILLER_0_106_192 ();
 sg13g2_fill_8 FILLER_0_106_200 ();
 sg13g2_fill_8 FILLER_0_106_208 ();
 sg13g2_fill_4 FILLER_0_106_216 ();
 sg13g2_fill_8 FILLER_0_106_225 ();
 sg13g2_fill_8 FILLER_0_106_233 ();
 sg13g2_fill_8 FILLER_0_106_241 ();
 sg13g2_fill_8 FILLER_0_106_249 ();
 sg13g2_fill_1 FILLER_0_106_257 ();
 sg13g2_fill_2 FILLER_0_106_263 ();
 sg13g2_fill_8 FILLER_0_106_269 ();
 sg13g2_fill_8 FILLER_0_106_277 ();
 sg13g2_fill_8 FILLER_0_106_285 ();
 sg13g2_fill_2 FILLER_0_106_298 ();
 sg13g2_fill_8 FILLER_0_106_326 ();
 sg13g2_fill_4 FILLER_0_106_334 ();
 sg13g2_fill_2 FILLER_0_106_338 ();
 sg13g2_fill_8 FILLER_0_106_345 ();
 sg13g2_fill_8 FILLER_0_106_353 ();
 sg13g2_fill_1 FILLER_0_106_361 ();
 sg13g2_fill_8 FILLER_0_106_366 ();
 sg13g2_fill_1 FILLER_0_106_374 ();
 sg13g2_fill_4 FILLER_0_106_380 ();
 sg13g2_fill_2 FILLER_0_106_384 ();
 sg13g2_fill_1 FILLER_0_106_386 ();
 sg13g2_fill_8 FILLER_0_106_392 ();
 sg13g2_fill_8 FILLER_0_106_400 ();
 sg13g2_fill_8 FILLER_0_106_408 ();
 sg13g2_fill_8 FILLER_0_106_420 ();
 sg13g2_fill_8 FILLER_0_106_428 ();
 sg13g2_fill_2 FILLER_0_106_441 ();
 sg13g2_fill_2 FILLER_0_106_447 ();
 sg13g2_fill_1 FILLER_0_106_449 ();
 sg13g2_fill_4 FILLER_0_106_476 ();
 sg13g2_fill_2 FILLER_0_106_480 ();
 sg13g2_fill_8 FILLER_0_106_485 ();
 sg13g2_fill_8 FILLER_0_106_493 ();
 sg13g2_fill_8 FILLER_0_106_501 ();
 sg13g2_fill_8 FILLER_0_106_509 ();
 sg13g2_fill_8 FILLER_0_106_517 ();
 sg13g2_fill_1 FILLER_0_106_525 ();
 sg13g2_fill_8 FILLER_0_106_530 ();
 sg13g2_fill_2 FILLER_0_106_543 ();
 sg13g2_fill_2 FILLER_0_106_549 ();
 sg13g2_fill_8 FILLER_0_106_557 ();
 sg13g2_fill_8 FILLER_0_106_565 ();
 sg13g2_fill_2 FILLER_0_106_573 ();
 sg13g2_fill_1 FILLER_0_106_575 ();
 sg13g2_fill_4 FILLER_0_106_580 ();
 sg13g2_fill_1 FILLER_0_106_584 ();
 sg13g2_fill_2 FILLER_0_106_589 ();
 sg13g2_fill_2 FILLER_0_106_617 ();
 sg13g2_fill_8 FILLER_0_106_624 ();
 sg13g2_fill_4 FILLER_0_106_632 ();
 sg13g2_fill_2 FILLER_0_106_636 ();
 sg13g2_fill_4 FILLER_0_106_664 ();
 sg13g2_fill_2 FILLER_0_106_668 ();
 sg13g2_fill_8 FILLER_0_106_675 ();
 sg13g2_fill_4 FILLER_0_106_683 ();
 sg13g2_fill_2 FILLER_0_106_693 ();
 sg13g2_fill_2 FILLER_0_106_721 ();
 sg13g2_fill_8 FILLER_0_106_728 ();
 sg13g2_fill_4 FILLER_0_106_741 ();
 sg13g2_fill_1 FILLER_0_106_745 ();
 sg13g2_fill_2 FILLER_0_106_750 ();
 sg13g2_fill_8 FILLER_0_106_758 ();
 sg13g2_fill_1 FILLER_0_106_766 ();
 sg13g2_fill_2 FILLER_0_106_771 ();
 sg13g2_fill_2 FILLER_0_106_778 ();
 sg13g2_fill_8 FILLER_0_106_785 ();
 sg13g2_fill_8 FILLER_0_106_793 ();
 sg13g2_fill_8 FILLER_0_106_801 ();
 sg13g2_fill_8 FILLER_0_106_809 ();
 sg13g2_fill_8 FILLER_0_106_817 ();
 sg13g2_fill_2 FILLER_0_106_825 ();
 sg13g2_fill_1 FILLER_0_106_827 ();
 sg13g2_fill_2 FILLER_0_106_833 ();
 sg13g2_fill_4 FILLER_0_106_839 ();
 sg13g2_fill_1 FILLER_0_106_843 ();
 sg13g2_fill_8 FILLER_0_106_849 ();
 sg13g2_fill_8 FILLER_0_106_857 ();
 sg13g2_fill_4 FILLER_0_106_865 ();
 sg13g2_fill_2 FILLER_0_106_869 ();
 sg13g2_fill_8 FILLER_0_106_877 ();
 sg13g2_fill_8 FILLER_0_106_885 ();
 sg13g2_fill_1 FILLER_0_106_893 ();
 sg13g2_fill_2 FILLER_0_106_898 ();
 sg13g2_fill_8 FILLER_0_106_905 ();
 sg13g2_fill_4 FILLER_0_106_913 ();
 sg13g2_fill_4 FILLER_0_106_922 ();
 sg13g2_fill_1 FILLER_0_106_926 ();
 sg13g2_fill_2 FILLER_0_106_937 ();
 sg13g2_fill_8 FILLER_0_106_949 ();
 sg13g2_fill_2 FILLER_0_106_957 ();
 sg13g2_fill_2 FILLER_0_106_963 ();
 sg13g2_fill_4 FILLER_0_106_969 ();
 sg13g2_fill_2 FILLER_0_106_983 ();
 sg13g2_fill_2 FILLER_0_106_989 ();
 sg13g2_fill_2 FILLER_0_106_995 ();
 sg13g2_fill_4 FILLER_0_106_1002 ();
 sg13g2_fill_2 FILLER_0_106_1014 ();
 sg13g2_fill_2 FILLER_0_106_1021 ();
 sg13g2_fill_1 FILLER_0_106_1023 ();
 sg13g2_fill_8 FILLER_0_106_1028 ();
 sg13g2_fill_2 FILLER_0_106_1036 ();
 sg13g2_fill_1 FILLER_0_106_1038 ();
 sg13g2_fill_2 FILLER_0_106_1045 ();
 sg13g2_fill_8 FILLER_0_106_1051 ();
 sg13g2_fill_4 FILLER_0_106_1059 ();
 sg13g2_fill_1 FILLER_0_106_1063 ();
 sg13g2_fill_2 FILLER_0_106_1069 ();
 sg13g2_fill_8 FILLER_0_106_1076 ();
 sg13g2_fill_2 FILLER_0_106_1088 ();
 sg13g2_fill_8 FILLER_0_106_1095 ();
 sg13g2_fill_8 FILLER_0_106_1103 ();
 sg13g2_fill_4 FILLER_0_106_1111 ();
 sg13g2_fill_2 FILLER_0_106_1115 ();
 sg13g2_fill_1 FILLER_0_106_1117 ();
 sg13g2_fill_8 FILLER_0_106_1125 ();
 sg13g2_fill_1 FILLER_0_106_1133 ();
 sg13g2_fill_8 FILLER_0_106_1139 ();
 sg13g2_fill_1 FILLER_0_106_1147 ();
 sg13g2_fill_8 FILLER_0_106_1153 ();
 sg13g2_fill_1 FILLER_0_106_1161 ();
 sg13g2_fill_8 FILLER_0_106_1170 ();
 sg13g2_fill_2 FILLER_0_106_1184 ();
 sg13g2_fill_8 FILLER_0_106_1190 ();
 sg13g2_fill_8 FILLER_0_106_1198 ();
 sg13g2_fill_8 FILLER_0_106_1206 ();
 sg13g2_fill_1 FILLER_0_106_1214 ();
 sg13g2_fill_2 FILLER_0_106_1222 ();
 sg13g2_fill_1 FILLER_0_106_1224 ();
 sg13g2_fill_2 FILLER_0_106_1231 ();
 sg13g2_fill_1 FILLER_0_106_1233 ();
 sg13g2_fill_2 FILLER_0_106_1240 ();
 sg13g2_fill_1 FILLER_0_106_1242 ();
 sg13g2_fill_2 FILLER_0_106_1251 ();
 sg13g2_fill_4 FILLER_0_106_1279 ();
 sg13g2_fill_8 FILLER_0_106_1287 ();
 sg13g2_fill_2 FILLER_0_106_1295 ();
 sg13g2_fill_8 FILLER_0_107_0 ();
 sg13g2_fill_8 FILLER_0_107_8 ();
 sg13g2_fill_8 FILLER_0_107_16 ();
 sg13g2_fill_8 FILLER_0_107_24 ();
 sg13g2_fill_8 FILLER_0_107_32 ();
 sg13g2_fill_8 FILLER_0_107_40 ();
 sg13g2_fill_8 FILLER_0_107_48 ();
 sg13g2_fill_8 FILLER_0_107_56 ();
 sg13g2_fill_8 FILLER_0_107_64 ();
 sg13g2_fill_8 FILLER_0_107_72 ();
 sg13g2_fill_8 FILLER_0_107_80 ();
 sg13g2_fill_8 FILLER_0_107_88 ();
 sg13g2_fill_8 FILLER_0_107_96 ();
 sg13g2_fill_8 FILLER_0_107_104 ();
 sg13g2_fill_8 FILLER_0_107_112 ();
 sg13g2_fill_8 FILLER_0_107_120 ();
 sg13g2_fill_8 FILLER_0_107_128 ();
 sg13g2_fill_8 FILLER_0_107_136 ();
 sg13g2_fill_8 FILLER_0_107_144 ();
 sg13g2_fill_8 FILLER_0_107_152 ();
 sg13g2_fill_8 FILLER_0_107_160 ();
 sg13g2_fill_8 FILLER_0_107_168 ();
 sg13g2_fill_8 FILLER_0_107_176 ();
 sg13g2_fill_8 FILLER_0_107_184 ();
 sg13g2_fill_8 FILLER_0_107_192 ();
 sg13g2_fill_8 FILLER_0_107_200 ();
 sg13g2_fill_2 FILLER_0_107_208 ();
 sg13g2_fill_2 FILLER_0_107_236 ();
 sg13g2_fill_8 FILLER_0_107_264 ();
 sg13g2_fill_8 FILLER_0_107_272 ();
 sg13g2_fill_8 FILLER_0_107_280 ();
 sg13g2_fill_8 FILLER_0_107_288 ();
 sg13g2_fill_8 FILLER_0_107_296 ();
 sg13g2_fill_2 FILLER_0_107_304 ();
 sg13g2_fill_1 FILLER_0_107_306 ();
 sg13g2_fill_8 FILLER_0_107_312 ();
 sg13g2_fill_8 FILLER_0_107_320 ();
 sg13g2_fill_8 FILLER_0_107_328 ();
 sg13g2_fill_4 FILLER_0_107_336 ();
 sg13g2_fill_1 FILLER_0_107_340 ();
 sg13g2_fill_8 FILLER_0_107_345 ();
 sg13g2_fill_8 FILLER_0_107_353 ();
 sg13g2_fill_8 FILLER_0_107_361 ();
 sg13g2_fill_8 FILLER_0_107_369 ();
 sg13g2_fill_2 FILLER_0_107_377 ();
 sg13g2_fill_2 FILLER_0_107_405 ();
 sg13g2_fill_8 FILLER_0_107_412 ();
 sg13g2_fill_8 FILLER_0_107_420 ();
 sg13g2_fill_8 FILLER_0_107_428 ();
 sg13g2_fill_4 FILLER_0_107_436 ();
 sg13g2_fill_1 FILLER_0_107_440 ();
 sg13g2_fill_2 FILLER_0_107_446 ();
 sg13g2_fill_4 FILLER_0_107_453 ();
 sg13g2_fill_8 FILLER_0_107_461 ();
 sg13g2_fill_2 FILLER_0_107_469 ();
 sg13g2_fill_8 FILLER_0_107_476 ();
 sg13g2_fill_1 FILLER_0_107_484 ();
 sg13g2_fill_8 FILLER_0_107_511 ();
 sg13g2_fill_8 FILLER_0_107_519 ();
 sg13g2_fill_8 FILLER_0_107_527 ();
 sg13g2_fill_8 FILLER_0_107_535 ();
 sg13g2_fill_8 FILLER_0_107_543 ();
 sg13g2_fill_8 FILLER_0_107_551 ();
 sg13g2_fill_8 FILLER_0_107_559 ();
 sg13g2_fill_8 FILLER_0_107_567 ();
 sg13g2_fill_2 FILLER_0_107_575 ();
 sg13g2_fill_8 FILLER_0_107_581 ();
 sg13g2_fill_8 FILLER_0_107_589 ();
 sg13g2_fill_8 FILLER_0_107_597 ();
 sg13g2_fill_8 FILLER_0_107_605 ();
 sg13g2_fill_8 FILLER_0_107_613 ();
 sg13g2_fill_8 FILLER_0_107_621 ();
 sg13g2_fill_4 FILLER_0_107_629 ();
 sg13g2_fill_1 FILLER_0_107_633 ();
 sg13g2_fill_4 FILLER_0_107_639 ();
 sg13g2_fill_2 FILLER_0_107_643 ();
 sg13g2_fill_4 FILLER_0_107_650 ();
 sg13g2_fill_2 FILLER_0_107_654 ();
 sg13g2_fill_8 FILLER_0_107_682 ();
 sg13g2_fill_4 FILLER_0_107_690 ();
 sg13g2_fill_2 FILLER_0_107_694 ();
 sg13g2_fill_1 FILLER_0_107_696 ();
 sg13g2_fill_2 FILLER_0_107_702 ();
 sg13g2_fill_8 FILLER_0_107_708 ();
 sg13g2_fill_8 FILLER_0_107_716 ();
 sg13g2_fill_2 FILLER_0_107_724 ();
 sg13g2_fill_1 FILLER_0_107_726 ();
 sg13g2_fill_2 FILLER_0_107_732 ();
 sg13g2_fill_2 FILLER_0_107_738 ();
 sg13g2_fill_8 FILLER_0_107_745 ();
 sg13g2_fill_1 FILLER_0_107_753 ();
 sg13g2_fill_8 FILLER_0_107_759 ();
 sg13g2_fill_4 FILLER_0_107_767 ();
 sg13g2_fill_2 FILLER_0_107_778 ();
 sg13g2_fill_1 FILLER_0_107_780 ();
 sg13g2_fill_2 FILLER_0_107_786 ();
 sg13g2_fill_1 FILLER_0_107_788 ();
 sg13g2_fill_2 FILLER_0_107_795 ();
 sg13g2_fill_1 FILLER_0_107_797 ();
 sg13g2_fill_2 FILLER_0_107_819 ();
 sg13g2_fill_2 FILLER_0_107_847 ();
 sg13g2_fill_8 FILLER_0_107_854 ();
 sg13g2_fill_2 FILLER_0_107_869 ();
 sg13g2_fill_8 FILLER_0_107_876 ();
 sg13g2_fill_4 FILLER_0_107_884 ();
 sg13g2_fill_4 FILLER_0_107_892 ();
 sg13g2_fill_8 FILLER_0_107_901 ();
 sg13g2_fill_2 FILLER_0_107_930 ();
 sg13g2_fill_4 FILLER_0_107_937 ();
 sg13g2_fill_8 FILLER_0_107_946 ();
 sg13g2_fill_4 FILLER_0_107_954 ();
 sg13g2_fill_2 FILLER_0_107_963 ();
 sg13g2_fill_2 FILLER_0_107_971 ();
 sg13g2_fill_1 FILLER_0_107_973 ();
 sg13g2_fill_2 FILLER_0_107_979 ();
 sg13g2_fill_2 FILLER_0_107_985 ();
 sg13g2_fill_8 FILLER_0_107_991 ();
 sg13g2_fill_4 FILLER_0_107_999 ();
 sg13g2_fill_8 FILLER_0_107_1008 ();
 sg13g2_fill_8 FILLER_0_107_1016 ();
 sg13g2_fill_8 FILLER_0_107_1024 ();
 sg13g2_fill_8 FILLER_0_107_1032 ();
 sg13g2_fill_8 FILLER_0_107_1040 ();
 sg13g2_fill_8 FILLER_0_107_1048 ();
 sg13g2_fill_8 FILLER_0_107_1056 ();
 sg13g2_fill_2 FILLER_0_107_1068 ();
 sg13g2_fill_2 FILLER_0_107_1078 ();
 sg13g2_fill_4 FILLER_0_107_1085 ();
 sg13g2_fill_2 FILLER_0_107_1089 ();
 sg13g2_fill_1 FILLER_0_107_1091 ();
 sg13g2_fill_8 FILLER_0_107_1096 ();
 sg13g2_fill_8 FILLER_0_107_1104 ();
 sg13g2_fill_1 FILLER_0_107_1112 ();
 sg13g2_fill_2 FILLER_0_107_1118 ();
 sg13g2_fill_1 FILLER_0_107_1120 ();
 sg13g2_fill_2 FILLER_0_107_1126 ();
 sg13g2_fill_2 FILLER_0_107_1135 ();
 sg13g2_fill_8 FILLER_0_107_1144 ();
 sg13g2_fill_8 FILLER_0_107_1152 ();
 sg13g2_fill_8 FILLER_0_107_1160 ();
 sg13g2_fill_8 FILLER_0_107_1168 ();
 sg13g2_fill_4 FILLER_0_107_1176 ();
 sg13g2_fill_1 FILLER_0_107_1180 ();
 sg13g2_fill_8 FILLER_0_107_1185 ();
 sg13g2_fill_8 FILLER_0_107_1193 ();
 sg13g2_fill_8 FILLER_0_107_1201 ();
 sg13g2_fill_8 FILLER_0_107_1209 ();
 sg13g2_fill_8 FILLER_0_107_1217 ();
 sg13g2_fill_2 FILLER_0_107_1225 ();
 sg13g2_fill_2 FILLER_0_107_1233 ();
 sg13g2_fill_2 FILLER_0_107_1240 ();
 sg13g2_fill_4 FILLER_0_107_1247 ();
 sg13g2_fill_1 FILLER_0_107_1251 ();
 sg13g2_fill_2 FILLER_0_107_1262 ();
 sg13g2_fill_2 FILLER_0_107_1268 ();
 sg13g2_fill_1 FILLER_0_107_1270 ();
 sg13g2_fill_2 FILLER_0_107_1275 ();
 sg13g2_fill_1 FILLER_0_107_1277 ();
 sg13g2_fill_2 FILLER_0_107_1282 ();
 sg13g2_fill_2 FILLER_0_107_1288 ();
 sg13g2_fill_2 FILLER_0_107_1294 ();
 sg13g2_fill_1 FILLER_0_107_1296 ();
 sg13g2_fill_8 FILLER_0_108_0 ();
 sg13g2_fill_8 FILLER_0_108_8 ();
 sg13g2_fill_8 FILLER_0_108_16 ();
 sg13g2_fill_8 FILLER_0_108_24 ();
 sg13g2_fill_8 FILLER_0_108_32 ();
 sg13g2_fill_8 FILLER_0_108_40 ();
 sg13g2_fill_8 FILLER_0_108_48 ();
 sg13g2_fill_8 FILLER_0_108_56 ();
 sg13g2_fill_8 FILLER_0_108_64 ();
 sg13g2_fill_8 FILLER_0_108_72 ();
 sg13g2_fill_8 FILLER_0_108_80 ();
 sg13g2_fill_8 FILLER_0_108_88 ();
 sg13g2_fill_8 FILLER_0_108_96 ();
 sg13g2_fill_8 FILLER_0_108_104 ();
 sg13g2_fill_8 FILLER_0_108_112 ();
 sg13g2_fill_8 FILLER_0_108_120 ();
 sg13g2_fill_8 FILLER_0_108_128 ();
 sg13g2_fill_8 FILLER_0_108_136 ();
 sg13g2_fill_8 FILLER_0_108_144 ();
 sg13g2_fill_8 FILLER_0_108_152 ();
 sg13g2_fill_8 FILLER_0_108_160 ();
 sg13g2_fill_8 FILLER_0_108_168 ();
 sg13g2_fill_8 FILLER_0_108_176 ();
 sg13g2_fill_8 FILLER_0_108_184 ();
 sg13g2_fill_8 FILLER_0_108_192 ();
 sg13g2_fill_8 FILLER_0_108_200 ();
 sg13g2_fill_8 FILLER_0_108_208 ();
 sg13g2_fill_8 FILLER_0_108_216 ();
 sg13g2_fill_8 FILLER_0_108_228 ();
 sg13g2_fill_2 FILLER_0_108_236 ();
 sg13g2_fill_1 FILLER_0_108_238 ();
 sg13g2_fill_2 FILLER_0_108_244 ();
 sg13g2_fill_1 FILLER_0_108_246 ();
 sg13g2_fill_2 FILLER_0_108_253 ();
 sg13g2_fill_1 FILLER_0_108_255 ();
 sg13g2_fill_2 FILLER_0_108_282 ();
 sg13g2_fill_4 FILLER_0_108_294 ();
 sg13g2_fill_4 FILLER_0_108_303 ();
 sg13g2_fill_8 FILLER_0_108_313 ();
 sg13g2_fill_8 FILLER_0_108_321 ();
 sg13g2_fill_8 FILLER_0_108_329 ();
 sg13g2_fill_8 FILLER_0_108_337 ();
 sg13g2_fill_8 FILLER_0_108_345 ();
 sg13g2_fill_8 FILLER_0_108_353 ();
 sg13g2_fill_8 FILLER_0_108_361 ();
 sg13g2_fill_8 FILLER_0_108_369 ();
 sg13g2_fill_8 FILLER_0_108_377 ();
 sg13g2_fill_2 FILLER_0_108_385 ();
 sg13g2_fill_8 FILLER_0_108_413 ();
 sg13g2_fill_2 FILLER_0_108_426 ();
 sg13g2_fill_2 FILLER_0_108_454 ();
 sg13g2_fill_2 FILLER_0_108_460 ();
 sg13g2_fill_2 FILLER_0_108_467 ();
 sg13g2_fill_8 FILLER_0_108_473 ();
 sg13g2_fill_8 FILLER_0_108_486 ();
 sg13g2_fill_8 FILLER_0_108_494 ();
 sg13g2_fill_8 FILLER_0_108_502 ();
 sg13g2_fill_8 FILLER_0_108_520 ();
 sg13g2_fill_8 FILLER_0_108_528 ();
 sg13g2_fill_4 FILLER_0_108_536 ();
 sg13g2_fill_2 FILLER_0_108_545 ();
 sg13g2_fill_8 FILLER_0_108_551 ();
 sg13g2_fill_2 FILLER_0_108_559 ();
 sg13g2_fill_1 FILLER_0_108_561 ();
 sg13g2_fill_8 FILLER_0_108_567 ();
 sg13g2_fill_8 FILLER_0_108_575 ();
 sg13g2_fill_1 FILLER_0_108_583 ();
 sg13g2_fill_8 FILLER_0_108_589 ();
 sg13g2_fill_8 FILLER_0_108_597 ();
 sg13g2_fill_4 FILLER_0_108_605 ();
 sg13g2_fill_2 FILLER_0_108_614 ();
 sg13g2_fill_2 FILLER_0_108_642 ();
 sg13g2_fill_2 FILLER_0_108_648 ();
 sg13g2_fill_8 FILLER_0_108_671 ();
 sg13g2_fill_8 FILLER_0_108_679 ();
 sg13g2_fill_8 FILLER_0_108_687 ();
 sg13g2_fill_4 FILLER_0_108_695 ();
 sg13g2_fill_4 FILLER_0_108_720 ();
 sg13g2_fill_8 FILLER_0_108_750 ();
 sg13g2_fill_8 FILLER_0_108_758 ();
 sg13g2_fill_8 FILLER_0_108_766 ();
 sg13g2_fill_8 FILLER_0_108_774 ();
 sg13g2_fill_2 FILLER_0_108_787 ();
 sg13g2_fill_8 FILLER_0_108_815 ();
 sg13g2_fill_2 FILLER_0_108_849 ();
 sg13g2_fill_8 FILLER_0_108_856 ();
 sg13g2_fill_8 FILLER_0_108_864 ();
 sg13g2_fill_8 FILLER_0_108_872 ();
 sg13g2_fill_8 FILLER_0_108_880 ();
 sg13g2_fill_2 FILLER_0_108_888 ();
 sg13g2_fill_2 FILLER_0_108_895 ();
 sg13g2_fill_2 FILLER_0_108_907 ();
 sg13g2_fill_4 FILLER_0_108_914 ();
 sg13g2_fill_1 FILLER_0_108_918 ();
 sg13g2_fill_4 FILLER_0_108_927 ();
 sg13g2_fill_2 FILLER_0_108_931 ();
 sg13g2_fill_1 FILLER_0_108_933 ();
 sg13g2_fill_2 FILLER_0_108_955 ();
 sg13g2_fill_1 FILLER_0_108_957 ();
 sg13g2_fill_2 FILLER_0_108_963 ();
 sg13g2_fill_8 FILLER_0_108_986 ();
 sg13g2_fill_2 FILLER_0_108_994 ();
 sg13g2_fill_2 FILLER_0_108_1000 ();
 sg13g2_fill_2 FILLER_0_108_1007 ();
 sg13g2_fill_2 FILLER_0_108_1014 ();
 sg13g2_fill_1 FILLER_0_108_1016 ();
 sg13g2_fill_8 FILLER_0_108_1022 ();
 sg13g2_fill_8 FILLER_0_108_1030 ();
 sg13g2_fill_8 FILLER_0_108_1038 ();
 sg13g2_fill_8 FILLER_0_108_1046 ();
 sg13g2_fill_8 FILLER_0_108_1054 ();
 sg13g2_fill_4 FILLER_0_108_1062 ();
 sg13g2_fill_1 FILLER_0_108_1066 ();
 sg13g2_fill_2 FILLER_0_108_1075 ();
 sg13g2_fill_8 FILLER_0_108_1081 ();
 sg13g2_fill_2 FILLER_0_108_1089 ();
 sg13g2_fill_2 FILLER_0_108_1096 ();
 sg13g2_fill_8 FILLER_0_108_1103 ();
 sg13g2_fill_8 FILLER_0_108_1111 ();
 sg13g2_fill_2 FILLER_0_108_1124 ();
 sg13g2_fill_8 FILLER_0_108_1133 ();
 sg13g2_fill_2 FILLER_0_108_1141 ();
 sg13g2_fill_4 FILLER_0_108_1147 ();
 sg13g2_fill_2 FILLER_0_108_1151 ();
 sg13g2_fill_1 FILLER_0_108_1153 ();
 sg13g2_fill_2 FILLER_0_108_1159 ();
 sg13g2_fill_8 FILLER_0_108_1166 ();
 sg13g2_fill_2 FILLER_0_108_1179 ();
 sg13g2_fill_4 FILLER_0_108_1186 ();
 sg13g2_fill_2 FILLER_0_108_1190 ();
 sg13g2_fill_1 FILLER_0_108_1192 ();
 sg13g2_fill_8 FILLER_0_108_1199 ();
 sg13g2_fill_4 FILLER_0_108_1207 ();
 sg13g2_fill_2 FILLER_0_108_1211 ();
 sg13g2_fill_8 FILLER_0_108_1218 ();
 sg13g2_fill_2 FILLER_0_108_1226 ();
 sg13g2_fill_2 FILLER_0_108_1234 ();
 sg13g2_fill_8 FILLER_0_108_1241 ();
 sg13g2_fill_2 FILLER_0_108_1249 ();
 sg13g2_fill_1 FILLER_0_108_1251 ();
 sg13g2_fill_2 FILLER_0_108_1262 ();
 sg13g2_fill_4 FILLER_0_108_1268 ();
 sg13g2_fill_2 FILLER_0_108_1272 ();
 sg13g2_fill_1 FILLER_0_108_1274 ();
 sg13g2_fill_8 FILLER_0_108_1283 ();
 sg13g2_fill_4 FILLER_0_108_1291 ();
 sg13g2_fill_2 FILLER_0_108_1295 ();
 sg13g2_fill_8 FILLER_0_109_0 ();
 sg13g2_fill_8 FILLER_0_109_8 ();
 sg13g2_fill_8 FILLER_0_109_16 ();
 sg13g2_fill_8 FILLER_0_109_24 ();
 sg13g2_fill_8 FILLER_0_109_32 ();
 sg13g2_fill_8 FILLER_0_109_40 ();
 sg13g2_fill_8 FILLER_0_109_48 ();
 sg13g2_fill_8 FILLER_0_109_56 ();
 sg13g2_fill_8 FILLER_0_109_64 ();
 sg13g2_fill_8 FILLER_0_109_72 ();
 sg13g2_fill_8 FILLER_0_109_80 ();
 sg13g2_fill_8 FILLER_0_109_88 ();
 sg13g2_fill_8 FILLER_0_109_96 ();
 sg13g2_fill_8 FILLER_0_109_104 ();
 sg13g2_fill_8 FILLER_0_109_112 ();
 sg13g2_fill_8 FILLER_0_109_120 ();
 sg13g2_fill_8 FILLER_0_109_128 ();
 sg13g2_fill_8 FILLER_0_109_136 ();
 sg13g2_fill_8 FILLER_0_109_144 ();
 sg13g2_fill_8 FILLER_0_109_152 ();
 sg13g2_fill_8 FILLER_0_109_160 ();
 sg13g2_fill_8 FILLER_0_109_168 ();
 sg13g2_fill_8 FILLER_0_109_176 ();
 sg13g2_fill_8 FILLER_0_109_184 ();
 sg13g2_fill_8 FILLER_0_109_192 ();
 sg13g2_fill_8 FILLER_0_109_200 ();
 sg13g2_fill_8 FILLER_0_109_208 ();
 sg13g2_fill_2 FILLER_0_109_216 ();
 sg13g2_fill_1 FILLER_0_109_218 ();
 sg13g2_fill_4 FILLER_0_109_245 ();
 sg13g2_fill_4 FILLER_0_109_270 ();
 sg13g2_fill_2 FILLER_0_109_279 ();
 sg13g2_fill_4 FILLER_0_109_285 ();
 sg13g2_fill_2 FILLER_0_109_295 ();
 sg13g2_fill_4 FILLER_0_109_303 ();
 sg13g2_fill_2 FILLER_0_109_307 ();
 sg13g2_fill_8 FILLER_0_109_314 ();
 sg13g2_fill_1 FILLER_0_109_322 ();
 sg13g2_fill_2 FILLER_0_109_328 ();
 sg13g2_fill_1 FILLER_0_109_330 ();
 sg13g2_fill_8 FILLER_0_109_335 ();
 sg13g2_fill_2 FILLER_0_109_343 ();
 sg13g2_fill_8 FILLER_0_109_350 ();
 sg13g2_fill_4 FILLER_0_109_358 ();
 sg13g2_fill_2 FILLER_0_109_362 ();
 sg13g2_fill_8 FILLER_0_109_368 ();
 sg13g2_fill_8 FILLER_0_109_376 ();
 sg13g2_fill_2 FILLER_0_109_389 ();
 sg13g2_fill_2 FILLER_0_109_396 ();
 sg13g2_fill_4 FILLER_0_109_402 ();
 sg13g2_fill_2 FILLER_0_109_406 ();
 sg13g2_fill_2 FILLER_0_109_412 ();
 sg13g2_fill_8 FILLER_0_109_424 ();
 sg13g2_fill_8 FILLER_0_109_432 ();
 sg13g2_fill_8 FILLER_0_109_440 ();
 sg13g2_fill_8 FILLER_0_109_448 ();
 sg13g2_fill_8 FILLER_0_109_456 ();
 sg13g2_fill_8 FILLER_0_109_464 ();
 sg13g2_fill_8 FILLER_0_109_472 ();
 sg13g2_fill_2 FILLER_0_109_480 ();
 sg13g2_fill_1 FILLER_0_109_482 ();
 sg13g2_fill_4 FILLER_0_109_488 ();
 sg13g2_fill_2 FILLER_0_109_492 ();
 sg13g2_fill_1 FILLER_0_109_494 ();
 sg13g2_fill_8 FILLER_0_109_521 ();
 sg13g2_fill_2 FILLER_0_109_529 ();
 sg13g2_fill_2 FILLER_0_109_536 ();
 sg13g2_fill_2 FILLER_0_109_564 ();
 sg13g2_fill_8 FILLER_0_109_576 ();
 sg13g2_fill_1 FILLER_0_109_584 ();
 sg13g2_fill_8 FILLER_0_109_611 ();
 sg13g2_fill_8 FILLER_0_109_619 ();
 sg13g2_fill_8 FILLER_0_109_627 ();
 sg13g2_fill_2 FILLER_0_109_639 ();
 sg13g2_fill_8 FILLER_0_109_645 ();
 sg13g2_fill_8 FILLER_0_109_653 ();
 sg13g2_fill_8 FILLER_0_109_661 ();
 sg13g2_fill_2 FILLER_0_109_669 ();
 sg13g2_fill_1 FILLER_0_109_671 ();
 sg13g2_fill_4 FILLER_0_109_677 ();
 sg13g2_fill_2 FILLER_0_109_686 ();
 sg13g2_fill_4 FILLER_0_109_692 ();
 sg13g2_fill_1 FILLER_0_109_696 ();
 sg13g2_fill_2 FILLER_0_109_702 ();
 sg13g2_fill_4 FILLER_0_109_709 ();
 sg13g2_fill_2 FILLER_0_109_713 ();
 sg13g2_fill_8 FILLER_0_109_725 ();
 sg13g2_fill_4 FILLER_0_109_733 ();
 sg13g2_fill_8 FILLER_0_109_742 ();
 sg13g2_fill_8 FILLER_0_109_750 ();
 sg13g2_fill_8 FILLER_0_109_758 ();
 sg13g2_fill_4 FILLER_0_109_766 ();
 sg13g2_fill_1 FILLER_0_109_770 ();
 sg13g2_fill_2 FILLER_0_109_776 ();
 sg13g2_fill_1 FILLER_0_109_778 ();
 sg13g2_fill_4 FILLER_0_109_805 ();
 sg13g2_fill_8 FILLER_0_109_813 ();
 sg13g2_fill_1 FILLER_0_109_821 ();
 sg13g2_fill_2 FILLER_0_109_827 ();
 sg13g2_fill_2 FILLER_0_109_834 ();
 sg13g2_fill_2 FILLER_0_109_841 ();
 sg13g2_fill_2 FILLER_0_109_847 ();
 sg13g2_fill_2 FILLER_0_109_853 ();
 sg13g2_fill_2 FILLER_0_109_860 ();
 sg13g2_fill_1 FILLER_0_109_862 ();
 sg13g2_fill_2 FILLER_0_109_867 ();
 sg13g2_fill_2 FILLER_0_109_874 ();
 sg13g2_fill_4 FILLER_0_109_880 ();
 sg13g2_fill_2 FILLER_0_109_884 ();
 sg13g2_fill_1 FILLER_0_109_886 ();
 sg13g2_fill_8 FILLER_0_109_891 ();
 sg13g2_fill_2 FILLER_0_109_899 ();
 sg13g2_fill_8 FILLER_0_109_906 ();
 sg13g2_fill_1 FILLER_0_109_914 ();
 sg13g2_fill_2 FILLER_0_109_920 ();
 sg13g2_fill_8 FILLER_0_109_943 ();
 sg13g2_fill_8 FILLER_0_109_951 ();
 sg13g2_fill_1 FILLER_0_109_959 ();
 sg13g2_fill_2 FILLER_0_109_966 ();
 sg13g2_fill_8 FILLER_0_109_972 ();
 sg13g2_fill_8 FILLER_0_109_980 ();
 sg13g2_fill_8 FILLER_0_109_988 ();
 sg13g2_fill_4 FILLER_0_109_996 ();
 sg13g2_fill_8 FILLER_0_109_1004 ();
 sg13g2_fill_2 FILLER_0_109_1020 ();
 sg13g2_fill_2 FILLER_0_109_1027 ();
 sg13g2_fill_8 FILLER_0_109_1035 ();
 sg13g2_fill_8 FILLER_0_109_1043 ();
 sg13g2_fill_8 FILLER_0_109_1051 ();
 sg13g2_fill_4 FILLER_0_109_1059 ();
 sg13g2_fill_2 FILLER_0_109_1063 ();
 sg13g2_fill_1 FILLER_0_109_1065 ();
 sg13g2_fill_2 FILLER_0_109_1074 ();
 sg13g2_fill_2 FILLER_0_109_1084 ();
 sg13g2_fill_4 FILLER_0_109_1091 ();
 sg13g2_fill_1 FILLER_0_109_1095 ();
 sg13g2_fill_4 FILLER_0_109_1102 ();
 sg13g2_fill_8 FILLER_0_109_1110 ();
 sg13g2_fill_8 FILLER_0_109_1118 ();
 sg13g2_fill_8 FILLER_0_109_1126 ();
 sg13g2_fill_8 FILLER_0_109_1134 ();
 sg13g2_fill_8 FILLER_0_109_1142 ();
 sg13g2_fill_8 FILLER_0_109_1150 ();
 sg13g2_fill_1 FILLER_0_109_1158 ();
 sg13g2_fill_8 FILLER_0_109_1165 ();
 sg13g2_fill_2 FILLER_0_109_1178 ();
 sg13g2_fill_2 FILLER_0_109_1188 ();
 sg13g2_fill_2 FILLER_0_109_1195 ();
 sg13g2_fill_1 FILLER_0_109_1197 ();
 sg13g2_fill_8 FILLER_0_109_1203 ();
 sg13g2_fill_8 FILLER_0_109_1211 ();
 sg13g2_fill_2 FILLER_0_109_1219 ();
 sg13g2_fill_2 FILLER_0_109_1226 ();
 sg13g2_fill_2 FILLER_0_109_1236 ();
 sg13g2_fill_8 FILLER_0_109_1243 ();
 sg13g2_fill_2 FILLER_0_109_1258 ();
 sg13g2_fill_2 FILLER_0_109_1265 ();
 sg13g2_fill_1 FILLER_0_109_1267 ();
 sg13g2_fill_4 FILLER_0_109_1273 ();
 sg13g2_fill_2 FILLER_0_109_1277 ();
 sg13g2_fill_4 FILLER_0_109_1285 ();
 sg13g2_fill_1 FILLER_0_109_1289 ();
 sg13g2_fill_2 FILLER_0_109_1294 ();
 sg13g2_fill_1 FILLER_0_109_1296 ();
 sg13g2_fill_8 FILLER_0_110_0 ();
 sg13g2_fill_8 FILLER_0_110_8 ();
 sg13g2_fill_8 FILLER_0_110_16 ();
 sg13g2_fill_8 FILLER_0_110_24 ();
 sg13g2_fill_8 FILLER_0_110_32 ();
 sg13g2_fill_8 FILLER_0_110_40 ();
 sg13g2_fill_8 FILLER_0_110_48 ();
 sg13g2_fill_8 FILLER_0_110_56 ();
 sg13g2_fill_8 FILLER_0_110_64 ();
 sg13g2_fill_8 FILLER_0_110_72 ();
 sg13g2_fill_8 FILLER_0_110_80 ();
 sg13g2_fill_8 FILLER_0_110_88 ();
 sg13g2_fill_8 FILLER_0_110_96 ();
 sg13g2_fill_8 FILLER_0_110_104 ();
 sg13g2_fill_8 FILLER_0_110_112 ();
 sg13g2_fill_8 FILLER_0_110_120 ();
 sg13g2_fill_8 FILLER_0_110_128 ();
 sg13g2_fill_8 FILLER_0_110_136 ();
 sg13g2_fill_8 FILLER_0_110_144 ();
 sg13g2_fill_8 FILLER_0_110_152 ();
 sg13g2_fill_8 FILLER_0_110_160 ();
 sg13g2_fill_8 FILLER_0_110_168 ();
 sg13g2_fill_8 FILLER_0_110_176 ();
 sg13g2_fill_8 FILLER_0_110_184 ();
 sg13g2_fill_8 FILLER_0_110_192 ();
 sg13g2_fill_8 FILLER_0_110_200 ();
 sg13g2_fill_8 FILLER_0_110_208 ();
 sg13g2_fill_8 FILLER_0_110_216 ();
 sg13g2_fill_2 FILLER_0_110_224 ();
 sg13g2_fill_2 FILLER_0_110_231 ();
 sg13g2_fill_8 FILLER_0_110_237 ();
 sg13g2_fill_8 FILLER_0_110_245 ();
 sg13g2_fill_8 FILLER_0_110_253 ();
 sg13g2_fill_8 FILLER_0_110_261 ();
 sg13g2_fill_8 FILLER_0_110_269 ();
 sg13g2_fill_1 FILLER_0_110_277 ();
 sg13g2_fill_2 FILLER_0_110_283 ();
 sg13g2_fill_4 FILLER_0_110_289 ();
 sg13g2_fill_1 FILLER_0_110_293 ();
 sg13g2_fill_2 FILLER_0_110_320 ();
 sg13g2_fill_2 FILLER_0_110_348 ();
 sg13g2_fill_4 FILLER_0_110_353 ();
 sg13g2_fill_2 FILLER_0_110_357 ();
 sg13g2_fill_4 FILLER_0_110_365 ();
 sg13g2_fill_2 FILLER_0_110_369 ();
 sg13g2_fill_8 FILLER_0_110_381 ();
 sg13g2_fill_8 FILLER_0_110_389 ();
 sg13g2_fill_2 FILLER_0_110_397 ();
 sg13g2_fill_1 FILLER_0_110_399 ();
 sg13g2_fill_8 FILLER_0_110_408 ();
 sg13g2_fill_4 FILLER_0_110_416 ();
 sg13g2_fill_2 FILLER_0_110_425 ();
 sg13g2_fill_8 FILLER_0_110_431 ();
 sg13g2_fill_8 FILLER_0_110_443 ();
 sg13g2_fill_8 FILLER_0_110_451 ();
 sg13g2_fill_8 FILLER_0_110_459 ();
 sg13g2_fill_8 FILLER_0_110_467 ();
 sg13g2_fill_8 FILLER_0_110_475 ();
 sg13g2_fill_8 FILLER_0_110_483 ();
 sg13g2_fill_8 FILLER_0_110_491 ();
 sg13g2_fill_8 FILLER_0_110_499 ();
 sg13g2_fill_2 FILLER_0_110_507 ();
 sg13g2_fill_1 FILLER_0_110_509 ();
 sg13g2_fill_4 FILLER_0_110_515 ();
 sg13g2_fill_2 FILLER_0_110_519 ();
 sg13g2_fill_2 FILLER_0_110_547 ();
 sg13g2_fill_8 FILLER_0_110_570 ();
 sg13g2_fill_2 FILLER_0_110_578 ();
 sg13g2_fill_1 FILLER_0_110_580 ();
 sg13g2_fill_4 FILLER_0_110_586 ();
 sg13g2_fill_2 FILLER_0_110_590 ();
 sg13g2_fill_2 FILLER_0_110_597 ();
 sg13g2_fill_1 FILLER_0_110_599 ();
 sg13g2_fill_2 FILLER_0_110_604 ();
 sg13g2_fill_1 FILLER_0_110_606 ();
 sg13g2_fill_8 FILLER_0_110_611 ();
 sg13g2_fill_4 FILLER_0_110_619 ();
 sg13g2_fill_2 FILLER_0_110_623 ();
 sg13g2_fill_1 FILLER_0_110_625 ();
 sg13g2_fill_8 FILLER_0_110_630 ();
 sg13g2_fill_2 FILLER_0_110_638 ();
 sg13g2_fill_1 FILLER_0_110_640 ();
 sg13g2_fill_2 FILLER_0_110_646 ();
 sg13g2_fill_1 FILLER_0_110_648 ();
 sg13g2_fill_8 FILLER_0_110_653 ();
 sg13g2_fill_8 FILLER_0_110_661 ();
 sg13g2_fill_8 FILLER_0_110_669 ();
 sg13g2_fill_2 FILLER_0_110_677 ();
 sg13g2_fill_2 FILLER_0_110_705 ();
 sg13g2_fill_1 FILLER_0_110_707 ();
 sg13g2_fill_8 FILLER_0_110_713 ();
 sg13g2_fill_8 FILLER_0_110_721 ();
 sg13g2_fill_8 FILLER_0_110_729 ();
 sg13g2_fill_8 FILLER_0_110_737 ();
 sg13g2_fill_4 FILLER_0_110_745 ();
 sg13g2_fill_1 FILLER_0_110_749 ();
 sg13g2_fill_4 FILLER_0_110_755 ();
 sg13g2_fill_1 FILLER_0_110_759 ();
 sg13g2_fill_8 FILLER_0_110_764 ();
 sg13g2_fill_8 FILLER_0_110_772 ();
 sg13g2_fill_4 FILLER_0_110_780 ();
 sg13g2_fill_2 FILLER_0_110_784 ();
 sg13g2_fill_1 FILLER_0_110_786 ();
 sg13g2_fill_4 FILLER_0_110_792 ();
 sg13g2_fill_4 FILLER_0_110_800 ();
 sg13g2_fill_2 FILLER_0_110_804 ();
 sg13g2_fill_1 FILLER_0_110_806 ();
 sg13g2_fill_2 FILLER_0_110_812 ();
 sg13g2_fill_2 FILLER_0_110_824 ();
 sg13g2_fill_1 FILLER_0_110_826 ();
 sg13g2_fill_8 FILLER_0_110_832 ();
 sg13g2_fill_2 FILLER_0_110_840 ();
 sg13g2_fill_8 FILLER_0_110_848 ();
 sg13g2_fill_8 FILLER_0_110_856 ();
 sg13g2_fill_2 FILLER_0_110_864 ();
 sg13g2_fill_1 FILLER_0_110_866 ();
 sg13g2_fill_8 FILLER_0_110_893 ();
 sg13g2_fill_4 FILLER_0_110_901 ();
 sg13g2_fill_4 FILLER_0_110_910 ();
 sg13g2_fill_2 FILLER_0_110_914 ();
 sg13g2_fill_1 FILLER_0_110_916 ();
 sg13g2_fill_2 FILLER_0_110_938 ();
 sg13g2_fill_2 FILLER_0_110_945 ();
 sg13g2_fill_4 FILLER_0_110_952 ();
 sg13g2_fill_2 FILLER_0_110_956 ();
 sg13g2_fill_1 FILLER_0_110_958 ();
 sg13g2_fill_2 FILLER_0_110_965 ();
 sg13g2_fill_8 FILLER_0_110_971 ();
 sg13g2_fill_8 FILLER_0_110_979 ();
 sg13g2_fill_8 FILLER_0_110_987 ();
 sg13g2_fill_4 FILLER_0_110_995 ();
 sg13g2_fill_4 FILLER_0_110_1007 ();
 sg13g2_fill_2 FILLER_0_110_1015 ();
 sg13g2_fill_8 FILLER_0_110_1023 ();
 sg13g2_fill_2 FILLER_0_110_1031 ();
 sg13g2_fill_1 FILLER_0_110_1033 ();
 sg13g2_fill_2 FILLER_0_110_1038 ();
 sg13g2_fill_2 FILLER_0_110_1047 ();
 sg13g2_fill_8 FILLER_0_110_1054 ();
 sg13g2_fill_2 FILLER_0_110_1062 ();
 sg13g2_fill_2 FILLER_0_110_1068 ();
 sg13g2_fill_2 FILLER_0_110_1075 ();
 sg13g2_fill_2 FILLER_0_110_1082 ();
 sg13g2_fill_1 FILLER_0_110_1084 ();
 sg13g2_fill_8 FILLER_0_110_1089 ();
 sg13g2_fill_8 FILLER_0_110_1097 ();
 sg13g2_fill_8 FILLER_0_110_1105 ();
 sg13g2_fill_8 FILLER_0_110_1113 ();
 sg13g2_fill_8 FILLER_0_110_1125 ();
 sg13g2_fill_8 FILLER_0_110_1133 ();
 sg13g2_fill_4 FILLER_0_110_1141 ();
 sg13g2_fill_8 FILLER_0_110_1150 ();
 sg13g2_fill_2 FILLER_0_110_1158 ();
 sg13g2_fill_2 FILLER_0_110_1166 ();
 sg13g2_fill_4 FILLER_0_110_1174 ();
 sg13g2_fill_2 FILLER_0_110_1178 ();
 sg13g2_fill_4 FILLER_0_110_1185 ();
 sg13g2_fill_2 FILLER_0_110_1189 ();
 sg13g2_fill_2 FILLER_0_110_1197 ();
 sg13g2_fill_8 FILLER_0_110_1203 ();
 sg13g2_fill_8 FILLER_0_110_1211 ();
 sg13g2_fill_8 FILLER_0_110_1219 ();
 sg13g2_fill_8 FILLER_0_110_1227 ();
 sg13g2_fill_2 FILLER_0_110_1235 ();
 sg13g2_fill_1 FILLER_0_110_1237 ();
 sg13g2_fill_8 FILLER_0_110_1242 ();
 sg13g2_fill_2 FILLER_0_110_1250 ();
 sg13g2_fill_4 FILLER_0_110_1257 ();
 sg13g2_fill_2 FILLER_0_110_1266 ();
 sg13g2_fill_2 FILLER_0_110_1274 ();
 sg13g2_fill_1 FILLER_0_110_1276 ();
 sg13g2_fill_4 FILLER_0_110_1286 ();
 sg13g2_fill_2 FILLER_0_110_1294 ();
 sg13g2_fill_1 FILLER_0_110_1296 ();
 sg13g2_fill_8 FILLER_0_111_0 ();
 sg13g2_fill_8 FILLER_0_111_8 ();
 sg13g2_fill_8 FILLER_0_111_16 ();
 sg13g2_fill_8 FILLER_0_111_24 ();
 sg13g2_fill_8 FILLER_0_111_32 ();
 sg13g2_fill_8 FILLER_0_111_40 ();
 sg13g2_fill_8 FILLER_0_111_48 ();
 sg13g2_fill_8 FILLER_0_111_56 ();
 sg13g2_fill_8 FILLER_0_111_64 ();
 sg13g2_fill_8 FILLER_0_111_72 ();
 sg13g2_fill_8 FILLER_0_111_80 ();
 sg13g2_fill_8 FILLER_0_111_88 ();
 sg13g2_fill_8 FILLER_0_111_96 ();
 sg13g2_fill_8 FILLER_0_111_104 ();
 sg13g2_fill_8 FILLER_0_111_112 ();
 sg13g2_fill_8 FILLER_0_111_120 ();
 sg13g2_fill_8 FILLER_0_111_128 ();
 sg13g2_fill_8 FILLER_0_111_136 ();
 sg13g2_fill_8 FILLER_0_111_144 ();
 sg13g2_fill_8 FILLER_0_111_152 ();
 sg13g2_fill_8 FILLER_0_111_160 ();
 sg13g2_fill_8 FILLER_0_111_168 ();
 sg13g2_fill_8 FILLER_0_111_176 ();
 sg13g2_fill_8 FILLER_0_111_184 ();
 sg13g2_fill_8 FILLER_0_111_192 ();
 sg13g2_fill_8 FILLER_0_111_200 ();
 sg13g2_fill_8 FILLER_0_111_208 ();
 sg13g2_fill_8 FILLER_0_111_216 ();
 sg13g2_fill_8 FILLER_0_111_224 ();
 sg13g2_fill_8 FILLER_0_111_232 ();
 sg13g2_fill_8 FILLER_0_111_240 ();
 sg13g2_fill_8 FILLER_0_111_248 ();
 sg13g2_fill_8 FILLER_0_111_256 ();
 sg13g2_fill_8 FILLER_0_111_264 ();
 sg13g2_fill_4 FILLER_0_111_272 ();
 sg13g2_fill_2 FILLER_0_111_302 ();
 sg13g2_fill_4 FILLER_0_111_309 ();
 sg13g2_fill_2 FILLER_0_111_313 ();
 sg13g2_fill_1 FILLER_0_111_315 ();
 sg13g2_fill_8 FILLER_0_111_337 ();
 sg13g2_fill_8 FILLER_0_111_371 ();
 sg13g2_fill_8 FILLER_0_111_379 ();
 sg13g2_fill_8 FILLER_0_111_387 ();
 sg13g2_fill_2 FILLER_0_111_395 ();
 sg13g2_fill_2 FILLER_0_111_418 ();
 sg13g2_fill_4 FILLER_0_111_426 ();
 sg13g2_fill_2 FILLER_0_111_434 ();
 sg13g2_fill_1 FILLER_0_111_436 ();
 sg13g2_fill_2 FILLER_0_111_445 ();
 sg13g2_fill_8 FILLER_0_111_459 ();
 sg13g2_fill_4 FILLER_0_111_467 ();
 sg13g2_fill_8 FILLER_0_111_476 ();
 sg13g2_fill_8 FILLER_0_111_484 ();
 sg13g2_fill_8 FILLER_0_111_492 ();
 sg13g2_fill_8 FILLER_0_111_500 ();
 sg13g2_fill_4 FILLER_0_111_508 ();
 sg13g2_fill_8 FILLER_0_111_517 ();
 sg13g2_fill_8 FILLER_0_111_525 ();
 sg13g2_fill_4 FILLER_0_111_538 ();
 sg13g2_fill_2 FILLER_0_111_542 ();
 sg13g2_fill_1 FILLER_0_111_544 ();
 sg13g2_fill_4 FILLER_0_111_549 ();
 sg13g2_fill_1 FILLER_0_111_553 ();
 sg13g2_fill_2 FILLER_0_111_558 ();
 sg13g2_fill_4 FILLER_0_111_570 ();
 sg13g2_fill_1 FILLER_0_111_574 ();
 sg13g2_fill_8 FILLER_0_111_601 ();
 sg13g2_fill_8 FILLER_0_111_609 ();
 sg13g2_fill_8 FILLER_0_111_622 ();
 sg13g2_fill_2 FILLER_0_111_630 ();
 sg13g2_fill_1 FILLER_0_111_632 ();
 sg13g2_fill_2 FILLER_0_111_638 ();
 sg13g2_fill_8 FILLER_0_111_666 ();
 sg13g2_fill_8 FILLER_0_111_674 ();
 sg13g2_fill_8 FILLER_0_111_682 ();
 sg13g2_fill_8 FILLER_0_111_690 ();
 sg13g2_fill_1 FILLER_0_111_698 ();
 sg13g2_fill_8 FILLER_0_111_707 ();
 sg13g2_fill_8 FILLER_0_111_727 ();
 sg13g2_fill_4 FILLER_0_111_735 ();
 sg13g2_fill_2 FILLER_0_111_739 ();
 sg13g2_fill_2 FILLER_0_111_767 ();
 sg13g2_fill_2 FILLER_0_111_773 ();
 sg13g2_fill_1 FILLER_0_111_775 ();
 sg13g2_fill_8 FILLER_0_111_781 ();
 sg13g2_fill_8 FILLER_0_111_789 ();
 sg13g2_fill_8 FILLER_0_111_797 ();
 sg13g2_fill_1 FILLER_0_111_805 ();
 sg13g2_fill_2 FILLER_0_111_813 ();
 sg13g2_fill_8 FILLER_0_111_820 ();
 sg13g2_fill_4 FILLER_0_111_828 ();
 sg13g2_fill_1 FILLER_0_111_832 ();
 sg13g2_fill_2 FILLER_0_111_841 ();
 sg13g2_fill_8 FILLER_0_111_849 ();
 sg13g2_fill_4 FILLER_0_111_857 ();
 sg13g2_fill_2 FILLER_0_111_866 ();
 sg13g2_fill_1 FILLER_0_111_868 ();
 sg13g2_fill_4 FILLER_0_111_874 ();
 sg13g2_fill_2 FILLER_0_111_878 ();
 sg13g2_fill_4 FILLER_0_111_887 ();
 sg13g2_fill_8 FILLER_0_111_894 ();
 sg13g2_fill_8 FILLER_0_111_902 ();
 sg13g2_fill_8 FILLER_0_111_910 ();
 sg13g2_fill_8 FILLER_0_111_918 ();
 sg13g2_fill_8 FILLER_0_111_926 ();
 sg13g2_fill_8 FILLER_0_111_934 ();
 sg13g2_fill_8 FILLER_0_111_942 ();
 sg13g2_fill_1 FILLER_0_111_950 ();
 sg13g2_fill_2 FILLER_0_111_955 ();
 sg13g2_fill_4 FILLER_0_111_961 ();
 sg13g2_fill_8 FILLER_0_111_973 ();
 sg13g2_fill_8 FILLER_0_111_981 ();
 sg13g2_fill_8 FILLER_0_111_989 ();
 sg13g2_fill_8 FILLER_0_111_997 ();
 sg13g2_fill_2 FILLER_0_111_1005 ();
 sg13g2_fill_1 FILLER_0_111_1007 ();
 sg13g2_fill_2 FILLER_0_111_1016 ();
 sg13g2_fill_2 FILLER_0_111_1022 ();
 sg13g2_fill_2 FILLER_0_111_1028 ();
 sg13g2_fill_2 FILLER_0_111_1035 ();
 sg13g2_fill_8 FILLER_0_111_1042 ();
 sg13g2_fill_8 FILLER_0_111_1050 ();
 sg13g2_fill_8 FILLER_0_111_1058 ();
 sg13g2_fill_8 FILLER_0_111_1066 ();
 sg13g2_fill_8 FILLER_0_111_1074 ();
 sg13g2_fill_8 FILLER_0_111_1082 ();
 sg13g2_fill_8 FILLER_0_111_1090 ();
 sg13g2_fill_2 FILLER_0_111_1098 ();
 sg13g2_fill_1 FILLER_0_111_1100 ();
 sg13g2_fill_2 FILLER_0_111_1111 ();
 sg13g2_fill_2 FILLER_0_111_1117 ();
 sg13g2_fill_2 FILLER_0_111_1124 ();
 sg13g2_fill_2 FILLER_0_111_1130 ();
 sg13g2_fill_2 FILLER_0_111_1137 ();
 sg13g2_fill_2 FILLER_0_111_1149 ();
 sg13g2_fill_8 FILLER_0_111_1155 ();
 sg13g2_fill_8 FILLER_0_111_1163 ();
 sg13g2_fill_8 FILLER_0_111_1171 ();
 sg13g2_fill_8 FILLER_0_111_1179 ();
 sg13g2_fill_8 FILLER_0_111_1187 ();
 sg13g2_fill_4 FILLER_0_111_1195 ();
 sg13g2_fill_1 FILLER_0_111_1199 ();
 sg13g2_fill_8 FILLER_0_111_1205 ();
 sg13g2_fill_2 FILLER_0_111_1216 ();
 sg13g2_fill_2 FILLER_0_111_1222 ();
 sg13g2_fill_4 FILLER_0_111_1230 ();
 sg13g2_fill_2 FILLER_0_111_1234 ();
 sg13g2_fill_1 FILLER_0_111_1236 ();
 sg13g2_fill_8 FILLER_0_111_1242 ();
 sg13g2_fill_2 FILLER_0_111_1250 ();
 sg13g2_fill_1 FILLER_0_111_1252 ();
 sg13g2_fill_2 FILLER_0_111_1257 ();
 sg13g2_fill_8 FILLER_0_111_1263 ();
 sg13g2_fill_4 FILLER_0_111_1275 ();
 sg13g2_fill_2 FILLER_0_111_1284 ();
 sg13g2_fill_2 FILLER_0_111_1290 ();
 sg13g2_fill_1 FILLER_0_111_1296 ();
 sg13g2_fill_8 FILLER_0_112_0 ();
 sg13g2_fill_8 FILLER_0_112_8 ();
 sg13g2_fill_8 FILLER_0_112_16 ();
 sg13g2_fill_8 FILLER_0_112_24 ();
 sg13g2_fill_8 FILLER_0_112_36 ();
 sg13g2_fill_8 FILLER_0_112_44 ();
 sg13g2_fill_8 FILLER_0_112_52 ();
 sg13g2_fill_8 FILLER_0_112_60 ();
 sg13g2_fill_8 FILLER_0_112_68 ();
 sg13g2_fill_8 FILLER_0_112_76 ();
 sg13g2_fill_8 FILLER_0_112_84 ();
 sg13g2_fill_8 FILLER_0_112_92 ();
 sg13g2_fill_8 FILLER_0_112_100 ();
 sg13g2_fill_8 FILLER_0_112_108 ();
 sg13g2_fill_8 FILLER_0_112_116 ();
 sg13g2_fill_8 FILLER_0_112_124 ();
 sg13g2_fill_8 FILLER_0_112_132 ();
 sg13g2_fill_8 FILLER_0_112_140 ();
 sg13g2_fill_8 FILLER_0_112_148 ();
 sg13g2_fill_8 FILLER_0_112_156 ();
 sg13g2_fill_8 FILLER_0_112_164 ();
 sg13g2_fill_8 FILLER_0_112_172 ();
 sg13g2_fill_8 FILLER_0_112_180 ();
 sg13g2_fill_8 FILLER_0_112_188 ();
 sg13g2_fill_8 FILLER_0_112_196 ();
 sg13g2_fill_8 FILLER_0_112_204 ();
 sg13g2_fill_8 FILLER_0_112_212 ();
 sg13g2_fill_8 FILLER_0_112_220 ();
 sg13g2_fill_8 FILLER_0_112_228 ();
 sg13g2_fill_1 FILLER_0_112_236 ();
 sg13g2_fill_4 FILLER_0_112_242 ();
 sg13g2_fill_2 FILLER_0_112_246 ();
 sg13g2_fill_8 FILLER_0_112_252 ();
 sg13g2_fill_8 FILLER_0_112_260 ();
 sg13g2_fill_8 FILLER_0_112_268 ();
 sg13g2_fill_8 FILLER_0_112_276 ();
 sg13g2_fill_8 FILLER_0_112_284 ();
 sg13g2_fill_8 FILLER_0_112_292 ();
 sg13g2_fill_4 FILLER_0_112_300 ();
 sg13g2_fill_2 FILLER_0_112_304 ();
 sg13g2_fill_8 FILLER_0_112_310 ();
 sg13g2_fill_8 FILLER_0_112_318 ();
 sg13g2_fill_8 FILLER_0_112_326 ();
 sg13g2_fill_8 FILLER_0_112_334 ();
 sg13g2_fill_8 FILLER_0_112_342 ();
 sg13g2_fill_4 FILLER_0_112_350 ();
 sg13g2_fill_8 FILLER_0_112_360 ();
 sg13g2_fill_8 FILLER_0_112_368 ();
 sg13g2_fill_4 FILLER_0_112_376 ();
 sg13g2_fill_2 FILLER_0_112_380 ();
 sg13g2_fill_1 FILLER_0_112_382 ();
 sg13g2_fill_8 FILLER_0_112_409 ();
 sg13g2_fill_2 FILLER_0_112_417 ();
 sg13g2_fill_1 FILLER_0_112_419 ();
 sg13g2_fill_8 FILLER_0_112_425 ();
 sg13g2_fill_8 FILLER_0_112_433 ();
 sg13g2_fill_8 FILLER_0_112_441 ();
 sg13g2_fill_8 FILLER_0_112_449 ();
 sg13g2_fill_2 FILLER_0_112_462 ();
 sg13g2_fill_2 FILLER_0_112_469 ();
 sg13g2_fill_2 FILLER_0_112_492 ();
 sg13g2_fill_2 FILLER_0_112_497 ();
 sg13g2_fill_8 FILLER_0_112_503 ();
 sg13g2_fill_2 FILLER_0_112_511 ();
 sg13g2_fill_1 FILLER_0_112_513 ();
 sg13g2_fill_4 FILLER_0_112_519 ();
 sg13g2_fill_2 FILLER_0_112_528 ();
 sg13g2_fill_8 FILLER_0_112_534 ();
 sg13g2_fill_8 FILLER_0_112_542 ();
 sg13g2_fill_4 FILLER_0_112_550 ();
 sg13g2_fill_2 FILLER_0_112_554 ();
 sg13g2_fill_8 FILLER_0_112_561 ();
 sg13g2_fill_1 FILLER_0_112_569 ();
 sg13g2_fill_8 FILLER_0_112_574 ();
 sg13g2_fill_8 FILLER_0_112_586 ();
 sg13g2_fill_2 FILLER_0_112_615 ();
 sg13g2_fill_8 FILLER_0_112_621 ();
 sg13g2_fill_8 FILLER_0_112_629 ();
 sg13g2_fill_8 FILLER_0_112_637 ();
 sg13g2_fill_8 FILLER_0_112_645 ();
 sg13g2_fill_8 FILLER_0_112_653 ();
 sg13g2_fill_8 FILLER_0_112_661 ();
 sg13g2_fill_4 FILLER_0_112_669 ();
 sg13g2_fill_2 FILLER_0_112_673 ();
 sg13g2_fill_2 FILLER_0_112_679 ();
 sg13g2_fill_8 FILLER_0_112_686 ();
 sg13g2_fill_8 FILLER_0_112_700 ();
 sg13g2_fill_8 FILLER_0_112_708 ();
 sg13g2_fill_4 FILLER_0_112_716 ();
 sg13g2_fill_2 FILLER_0_112_720 ();
 sg13g2_fill_2 FILLER_0_112_727 ();
 sg13g2_fill_2 FILLER_0_112_733 ();
 sg13g2_fill_2 FILLER_0_112_740 ();
 sg13g2_fill_2 FILLER_0_112_768 ();
 sg13g2_fill_4 FILLER_0_112_780 ();
 sg13g2_fill_2 FILLER_0_112_784 ();
 sg13g2_fill_4 FILLER_0_112_793 ();
 sg13g2_fill_8 FILLER_0_112_805 ();
 sg13g2_fill_8 FILLER_0_112_813 ();
 sg13g2_fill_8 FILLER_0_112_821 ();
 sg13g2_fill_1 FILLER_0_112_829 ();
 sg13g2_fill_2 FILLER_0_112_835 ();
 sg13g2_fill_4 FILLER_0_112_841 ();
 sg13g2_fill_1 FILLER_0_112_845 ();
 sg13g2_fill_8 FILLER_0_112_852 ();
 sg13g2_fill_2 FILLER_0_112_860 ();
 sg13g2_fill_1 FILLER_0_112_862 ();
 sg13g2_fill_8 FILLER_0_112_869 ();
 sg13g2_fill_4 FILLER_0_112_886 ();
 sg13g2_fill_2 FILLER_0_112_890 ();
 sg13g2_fill_8 FILLER_0_112_897 ();
 sg13g2_fill_8 FILLER_0_112_905 ();
 sg13g2_fill_8 FILLER_0_112_913 ();
 sg13g2_fill_1 FILLER_0_112_921 ();
 sg13g2_fill_2 FILLER_0_112_926 ();
 sg13g2_fill_8 FILLER_0_112_933 ();
 sg13g2_fill_4 FILLER_0_112_941 ();
 sg13g2_fill_2 FILLER_0_112_945 ();
 sg13g2_fill_2 FILLER_0_112_951 ();
 sg13g2_fill_2 FILLER_0_112_958 ();
 sg13g2_fill_2 FILLER_0_112_966 ();
 sg13g2_fill_8 FILLER_0_112_973 ();
 sg13g2_fill_8 FILLER_0_112_981 ();
 sg13g2_fill_8 FILLER_0_112_989 ();
 sg13g2_fill_8 FILLER_0_112_997 ();
 sg13g2_fill_8 FILLER_0_112_1005 ();
 sg13g2_fill_4 FILLER_0_112_1013 ();
 sg13g2_fill_1 FILLER_0_112_1017 ();
 sg13g2_fill_4 FILLER_0_112_1022 ();
 sg13g2_fill_2 FILLER_0_112_1026 ();
 sg13g2_fill_2 FILLER_0_112_1033 ();
 sg13g2_fill_2 FILLER_0_112_1042 ();
 sg13g2_fill_8 FILLER_0_112_1050 ();
 sg13g2_fill_8 FILLER_0_112_1058 ();
 sg13g2_fill_8 FILLER_0_112_1066 ();
 sg13g2_fill_8 FILLER_0_112_1074 ();
 sg13g2_fill_8 FILLER_0_112_1082 ();
 sg13g2_fill_4 FILLER_0_112_1090 ();
 sg13g2_fill_2 FILLER_0_112_1094 ();
 sg13g2_fill_1 FILLER_0_112_1096 ();
 sg13g2_fill_8 FILLER_0_112_1102 ();
 sg13g2_fill_8 FILLER_0_112_1110 ();
 sg13g2_fill_2 FILLER_0_112_1122 ();
 sg13g2_fill_1 FILLER_0_112_1124 ();
 sg13g2_fill_4 FILLER_0_112_1130 ();
 sg13g2_fill_2 FILLER_0_112_1139 ();
 sg13g2_fill_1 FILLER_0_112_1141 ();
 sg13g2_fill_4 FILLER_0_112_1147 ();
 sg13g2_fill_2 FILLER_0_112_1151 ();
 sg13g2_fill_2 FILLER_0_112_1158 ();
 sg13g2_fill_8 FILLER_0_112_1166 ();
 sg13g2_fill_8 FILLER_0_112_1174 ();
 sg13g2_fill_8 FILLER_0_112_1182 ();
 sg13g2_fill_8 FILLER_0_112_1194 ();
 sg13g2_fill_8 FILLER_0_112_1202 ();
 sg13g2_fill_2 FILLER_0_112_1210 ();
 sg13g2_fill_1 FILLER_0_112_1212 ();
 sg13g2_fill_8 FILLER_0_112_1219 ();
 sg13g2_fill_8 FILLER_0_112_1227 ();
 sg13g2_fill_8 FILLER_0_112_1235 ();
 sg13g2_fill_4 FILLER_0_112_1243 ();
 sg13g2_fill_2 FILLER_0_112_1247 ();
 sg13g2_fill_4 FILLER_0_112_1253 ();
 sg13g2_fill_2 FILLER_0_112_1257 ();
 sg13g2_fill_1 FILLER_0_112_1259 ();
 sg13g2_fill_2 FILLER_0_112_1265 ();
 sg13g2_fill_2 FILLER_0_112_1271 ();
 sg13g2_fill_2 FILLER_0_112_1278 ();
 sg13g2_fill_8 FILLER_0_112_1284 ();
 sg13g2_fill_1 FILLER_0_112_1296 ();
 sg13g2_fill_8 FILLER_0_113_0 ();
 sg13g2_fill_8 FILLER_0_113_8 ();
 sg13g2_fill_8 FILLER_0_113_16 ();
 sg13g2_fill_8 FILLER_0_113_24 ();
 sg13g2_fill_8 FILLER_0_113_32 ();
 sg13g2_fill_8 FILLER_0_113_40 ();
 sg13g2_fill_8 FILLER_0_113_48 ();
 sg13g2_fill_8 FILLER_0_113_56 ();
 sg13g2_fill_8 FILLER_0_113_64 ();
 sg13g2_fill_8 FILLER_0_113_72 ();
 sg13g2_fill_8 FILLER_0_113_80 ();
 sg13g2_fill_8 FILLER_0_113_88 ();
 sg13g2_fill_8 FILLER_0_113_96 ();
 sg13g2_fill_8 FILLER_0_113_104 ();
 sg13g2_fill_8 FILLER_0_113_112 ();
 sg13g2_fill_8 FILLER_0_113_120 ();
 sg13g2_fill_8 FILLER_0_113_128 ();
 sg13g2_fill_8 FILLER_0_113_136 ();
 sg13g2_fill_8 FILLER_0_113_144 ();
 sg13g2_fill_8 FILLER_0_113_152 ();
 sg13g2_fill_8 FILLER_0_113_160 ();
 sg13g2_fill_8 FILLER_0_113_168 ();
 sg13g2_fill_8 FILLER_0_113_176 ();
 sg13g2_fill_8 FILLER_0_113_184 ();
 sg13g2_fill_8 FILLER_0_113_192 ();
 sg13g2_fill_8 FILLER_0_113_200 ();
 sg13g2_fill_8 FILLER_0_113_208 ();
 sg13g2_fill_2 FILLER_0_113_216 ();
 sg13g2_fill_1 FILLER_0_113_218 ();
 sg13g2_fill_2 FILLER_0_113_224 ();
 sg13g2_fill_4 FILLER_0_113_230 ();
 sg13g2_fill_2 FILLER_0_113_260 ();
 sg13g2_fill_4 FILLER_0_113_268 ();
 sg13g2_fill_1 FILLER_0_113_272 ();
 sg13g2_fill_2 FILLER_0_113_278 ();
 sg13g2_fill_8 FILLER_0_113_284 ();
 sg13g2_fill_8 FILLER_0_113_292 ();
 sg13g2_fill_8 FILLER_0_113_300 ();
 sg13g2_fill_2 FILLER_0_113_308 ();
 sg13g2_fill_1 FILLER_0_113_310 ();
 sg13g2_fill_2 FILLER_0_113_316 ();
 sg13g2_fill_8 FILLER_0_113_322 ();
 sg13g2_fill_4 FILLER_0_113_330 ();
 sg13g2_fill_1 FILLER_0_113_334 ();
 sg13g2_fill_8 FILLER_0_113_340 ();
 sg13g2_fill_8 FILLER_0_113_348 ();
 sg13g2_fill_8 FILLER_0_113_356 ();
 sg13g2_fill_8 FILLER_0_113_364 ();
 sg13g2_fill_4 FILLER_0_113_372 ();
 sg13g2_fill_2 FILLER_0_113_376 ();
 sg13g2_fill_2 FILLER_0_113_404 ();
 sg13g2_fill_4 FILLER_0_113_416 ();
 sg13g2_fill_2 FILLER_0_113_425 ();
 sg13g2_fill_2 FILLER_0_113_432 ();
 sg13g2_fill_1 FILLER_0_113_434 ();
 sg13g2_fill_2 FILLER_0_113_439 ();
 sg13g2_fill_2 FILLER_0_113_446 ();
 sg13g2_fill_2 FILLER_0_113_474 ();
 sg13g2_fill_2 FILLER_0_113_480 ();
 sg13g2_fill_1 FILLER_0_113_482 ();
 sg13g2_fill_4 FILLER_0_113_509 ();
 sg13g2_fill_8 FILLER_0_113_539 ();
 sg13g2_fill_8 FILLER_0_113_547 ();
 sg13g2_fill_2 FILLER_0_113_555 ();
 sg13g2_fill_1 FILLER_0_113_557 ();
 sg13g2_fill_8 FILLER_0_113_566 ();
 sg13g2_fill_8 FILLER_0_113_574 ();
 sg13g2_fill_8 FILLER_0_113_582 ();
 sg13g2_fill_8 FILLER_0_113_590 ();
 sg13g2_fill_8 FILLER_0_113_598 ();
 sg13g2_fill_8 FILLER_0_113_606 ();
 sg13g2_fill_8 FILLER_0_113_614 ();
 sg13g2_fill_8 FILLER_0_113_622 ();
 sg13g2_fill_2 FILLER_0_113_630 ();
 sg13g2_fill_2 FILLER_0_113_638 ();
 sg13g2_fill_4 FILLER_0_113_646 ();
 sg13g2_fill_1 FILLER_0_113_650 ();
 sg13g2_fill_2 FILLER_0_113_656 ();
 sg13g2_fill_4 FILLER_0_113_662 ();
 sg13g2_fill_2 FILLER_0_113_666 ();
 sg13g2_fill_4 FILLER_0_113_672 ();
 sg13g2_fill_2 FILLER_0_113_681 ();
 sg13g2_fill_2 FILLER_0_113_709 ();
 sg13g2_fill_1 FILLER_0_113_711 ();
 sg13g2_fill_2 FILLER_0_113_717 ();
 sg13g2_fill_2 FILLER_0_113_745 ();
 sg13g2_fill_4 FILLER_0_113_752 ();
 sg13g2_fill_1 FILLER_0_113_756 ();
 sg13g2_fill_8 FILLER_0_113_778 ();
 sg13g2_fill_8 FILLER_0_113_786 ();
 sg13g2_fill_2 FILLER_0_113_794 ();
 sg13g2_fill_2 FILLER_0_113_802 ();
 sg13g2_fill_4 FILLER_0_113_810 ();
 sg13g2_fill_2 FILLER_0_113_814 ();
 sg13g2_fill_4 FILLER_0_113_821 ();
 sg13g2_fill_2 FILLER_0_113_825 ();
 sg13g2_fill_1 FILLER_0_113_827 ();
 sg13g2_fill_2 FILLER_0_113_832 ();
 sg13g2_fill_1 FILLER_0_113_834 ();
 sg13g2_fill_8 FILLER_0_113_861 ();
 sg13g2_fill_8 FILLER_0_113_869 ();
 sg13g2_fill_2 FILLER_0_113_877 ();
 sg13g2_fill_1 FILLER_0_113_879 ();
 sg13g2_fill_2 FILLER_0_113_884 ();
 sg13g2_fill_8 FILLER_0_113_892 ();
 sg13g2_fill_8 FILLER_0_113_907 ();
 sg13g2_fill_8 FILLER_0_113_915 ();
 sg13g2_fill_2 FILLER_0_113_923 ();
 sg13g2_fill_1 FILLER_0_113_925 ();
 sg13g2_fill_8 FILLER_0_113_931 ();
 sg13g2_fill_8 FILLER_0_113_939 ();
 sg13g2_fill_2 FILLER_0_113_947 ();
 sg13g2_fill_1 FILLER_0_113_949 ();
 sg13g2_fill_2 FILLER_0_113_954 ();
 sg13g2_fill_2 FILLER_0_113_961 ();
 sg13g2_fill_4 FILLER_0_113_966 ();
 sg13g2_fill_1 FILLER_0_113_970 ();
 sg13g2_fill_8 FILLER_0_113_976 ();
 sg13g2_fill_2 FILLER_0_113_984 ();
 sg13g2_fill_1 FILLER_0_113_986 ();
 sg13g2_fill_2 FILLER_0_113_994 ();
 sg13g2_fill_2 FILLER_0_113_1000 ();
 sg13g2_fill_2 FILLER_0_113_1010 ();
 sg13g2_fill_8 FILLER_0_113_1020 ();
 sg13g2_fill_4 FILLER_0_113_1028 ();
 sg13g2_fill_2 FILLER_0_113_1032 ();
 sg13g2_fill_2 FILLER_0_113_1041 ();
 sg13g2_fill_8 FILLER_0_113_1048 ();
 sg13g2_fill_4 FILLER_0_113_1056 ();
 sg13g2_fill_2 FILLER_0_113_1060 ();
 sg13g2_fill_2 FILLER_0_113_1068 ();
 sg13g2_fill_1 FILLER_0_113_1070 ();
 sg13g2_fill_2 FILLER_0_113_1077 ();
 sg13g2_fill_1 FILLER_0_113_1079 ();
 sg13g2_fill_8 FILLER_0_113_1085 ();
 sg13g2_fill_4 FILLER_0_113_1093 ();
 sg13g2_fill_2 FILLER_0_113_1097 ();
 sg13g2_fill_1 FILLER_0_113_1099 ();
 sg13g2_fill_2 FILLER_0_113_1104 ();
 sg13g2_fill_8 FILLER_0_113_1111 ();
 sg13g2_fill_4 FILLER_0_113_1119 ();
 sg13g2_fill_2 FILLER_0_113_1123 ();
 sg13g2_fill_2 FILLER_0_113_1130 ();
 sg13g2_fill_1 FILLER_0_113_1132 ();
 sg13g2_fill_4 FILLER_0_113_1138 ();
 sg13g2_fill_2 FILLER_0_113_1142 ();
 sg13g2_fill_1 FILLER_0_113_1144 ();
 sg13g2_fill_2 FILLER_0_113_1155 ();
 sg13g2_fill_2 FILLER_0_113_1165 ();
 sg13g2_fill_1 FILLER_0_113_1167 ();
 sg13g2_fill_2 FILLER_0_113_1178 ();
 sg13g2_fill_2 FILLER_0_113_1184 ();
 sg13g2_fill_1 FILLER_0_113_1186 ();
 sg13g2_fill_2 FILLER_0_113_1195 ();
 sg13g2_fill_4 FILLER_0_113_1202 ();
 sg13g2_fill_1 FILLER_0_113_1206 ();
 sg13g2_fill_2 FILLER_0_113_1214 ();
 sg13g2_fill_1 FILLER_0_113_1216 ();
 sg13g2_fill_4 FILLER_0_113_1220 ();
 sg13g2_fill_2 FILLER_0_113_1230 ();
 sg13g2_fill_8 FILLER_0_113_1237 ();
 sg13g2_fill_2 FILLER_0_113_1245 ();
 sg13g2_fill_1 FILLER_0_113_1247 ();
 sg13g2_fill_2 FILLER_0_113_1256 ();
 sg13g2_fill_2 FILLER_0_113_1264 ();
 sg13g2_fill_2 FILLER_0_113_1271 ();
 sg13g2_fill_2 FILLER_0_113_1278 ();
 sg13g2_fill_2 FILLER_0_113_1284 ();
 sg13g2_fill_2 FILLER_0_113_1290 ();
 sg13g2_fill_1 FILLER_0_113_1296 ();
 sg13g2_fill_8 FILLER_0_114_0 ();
 sg13g2_fill_8 FILLER_0_114_8 ();
 sg13g2_fill_8 FILLER_0_114_16 ();
 sg13g2_fill_8 FILLER_0_114_24 ();
 sg13g2_fill_8 FILLER_0_114_32 ();
 sg13g2_fill_8 FILLER_0_114_40 ();
 sg13g2_fill_8 FILLER_0_114_48 ();
 sg13g2_fill_8 FILLER_0_114_56 ();
 sg13g2_fill_8 FILLER_0_114_64 ();
 sg13g2_fill_8 FILLER_0_114_72 ();
 sg13g2_fill_8 FILLER_0_114_80 ();
 sg13g2_fill_8 FILLER_0_114_88 ();
 sg13g2_fill_8 FILLER_0_114_96 ();
 sg13g2_fill_8 FILLER_0_114_104 ();
 sg13g2_fill_8 FILLER_0_114_112 ();
 sg13g2_fill_8 FILLER_0_114_120 ();
 sg13g2_fill_8 FILLER_0_114_128 ();
 sg13g2_fill_8 FILLER_0_114_136 ();
 sg13g2_fill_8 FILLER_0_114_144 ();
 sg13g2_fill_8 FILLER_0_114_152 ();
 sg13g2_fill_8 FILLER_0_114_160 ();
 sg13g2_fill_8 FILLER_0_114_168 ();
 sg13g2_fill_8 FILLER_0_114_176 ();
 sg13g2_fill_8 FILLER_0_114_184 ();
 sg13g2_fill_8 FILLER_0_114_192 ();
 sg13g2_fill_8 FILLER_0_114_200 ();
 sg13g2_fill_4 FILLER_0_114_208 ();
 sg13g2_fill_2 FILLER_0_114_212 ();
 sg13g2_fill_8 FILLER_0_114_240 ();
 sg13g2_fill_1 FILLER_0_114_248 ();
 sg13g2_fill_2 FILLER_0_114_254 ();
 sg13g2_fill_2 FILLER_0_114_261 ();
 sg13g2_fill_2 FILLER_0_114_289 ();
 sg13g2_fill_1 FILLER_0_114_291 ();
 sg13g2_fill_4 FILLER_0_114_300 ();
 sg13g2_fill_2 FILLER_0_114_330 ();
 sg13g2_fill_4 FILLER_0_114_337 ();
 sg13g2_fill_2 FILLER_0_114_351 ();
 sg13g2_fill_8 FILLER_0_114_358 ();
 sg13g2_fill_4 FILLER_0_114_366 ();
 sg13g2_fill_2 FILLER_0_114_370 ();
 sg13g2_fill_1 FILLER_0_114_372 ();
 sg13g2_fill_2 FILLER_0_114_378 ();
 sg13g2_fill_8 FILLER_0_114_385 ();
 sg13g2_fill_2 FILLER_0_114_393 ();
 sg13g2_fill_1 FILLER_0_114_395 ();
 sg13g2_fill_2 FILLER_0_114_400 ();
 sg13g2_fill_8 FILLER_0_114_406 ();
 sg13g2_fill_8 FILLER_0_114_414 ();
 sg13g2_fill_2 FILLER_0_114_422 ();
 sg13g2_fill_8 FILLER_0_114_450 ();
 sg13g2_fill_4 FILLER_0_114_458 ();
 sg13g2_fill_4 FILLER_0_114_468 ();
 sg13g2_fill_4 FILLER_0_114_477 ();
 sg13g2_fill_2 FILLER_0_114_481 ();
 sg13g2_fill_8 FILLER_0_114_488 ();
 sg13g2_fill_4 FILLER_0_114_496 ();
 sg13g2_fill_2 FILLER_0_114_500 ();
 sg13g2_fill_8 FILLER_0_114_507 ();
 sg13g2_fill_8 FILLER_0_114_515 ();
 sg13g2_fill_1 FILLER_0_114_523 ();
 sg13g2_fill_2 FILLER_0_114_528 ();
 sg13g2_fill_1 FILLER_0_114_530 ();
 sg13g2_fill_2 FILLER_0_114_535 ();
 sg13g2_fill_2 FILLER_0_114_542 ();
 sg13g2_fill_8 FILLER_0_114_570 ();
 sg13g2_fill_4 FILLER_0_114_604 ();
 sg13g2_fill_2 FILLER_0_114_608 ();
 sg13g2_fill_8 FILLER_0_114_615 ();
 sg13g2_fill_8 FILLER_0_114_623 ();
 sg13g2_fill_8 FILLER_0_114_631 ();
 sg13g2_fill_4 FILLER_0_114_639 ();
 sg13g2_fill_2 FILLER_0_114_643 ();
 sg13g2_fill_1 FILLER_0_114_645 ();
 sg13g2_fill_2 FILLER_0_114_672 ();
 sg13g2_fill_2 FILLER_0_114_679 ();
 sg13g2_fill_1 FILLER_0_114_681 ();
 sg13g2_fill_4 FILLER_0_114_687 ();
 sg13g2_fill_2 FILLER_0_114_691 ();
 sg13g2_fill_1 FILLER_0_114_693 ();
 sg13g2_fill_8 FILLER_0_114_699 ();
 sg13g2_fill_8 FILLER_0_114_707 ();
 sg13g2_fill_8 FILLER_0_114_715 ();
 sg13g2_fill_2 FILLER_0_114_723 ();
 sg13g2_fill_1 FILLER_0_114_725 ();
 sg13g2_fill_2 FILLER_0_114_752 ();
 sg13g2_fill_8 FILLER_0_114_759 ();
 sg13g2_fill_4 FILLER_0_114_767 ();
 sg13g2_fill_8 FILLER_0_114_776 ();
 sg13g2_fill_8 FILLER_0_114_784 ();
 sg13g2_fill_2 FILLER_0_114_792 ();
 sg13g2_fill_1 FILLER_0_114_794 ();
 sg13g2_fill_2 FILLER_0_114_800 ();
 sg13g2_fill_2 FILLER_0_114_812 ();
 sg13g2_fill_2 FILLER_0_114_822 ();
 sg13g2_fill_2 FILLER_0_114_829 ();
 sg13g2_fill_8 FILLER_0_114_857 ();
 sg13g2_fill_1 FILLER_0_114_865 ();
 sg13g2_fill_2 FILLER_0_114_871 ();
 sg13g2_fill_2 FILLER_0_114_877 ();
 sg13g2_fill_2 FILLER_0_114_885 ();
 sg13g2_fill_1 FILLER_0_114_887 ();
 sg13g2_fill_8 FILLER_0_114_914 ();
 sg13g2_fill_4 FILLER_0_114_922 ();
 sg13g2_fill_4 FILLER_0_114_931 ();
 sg13g2_fill_1 FILLER_0_114_935 ();
 sg13g2_fill_2 FILLER_0_114_941 ();
 sg13g2_fill_8 FILLER_0_114_949 ();
 sg13g2_fill_4 FILLER_0_114_957 ();
 sg13g2_fill_2 FILLER_0_114_966 ();
 sg13g2_fill_2 FILLER_0_114_973 ();
 sg13g2_fill_8 FILLER_0_114_980 ();
 sg13g2_fill_4 FILLER_0_114_988 ();
 sg13g2_fill_2 FILLER_0_114_992 ();
 sg13g2_fill_1 FILLER_0_114_994 ();
 sg13g2_fill_2 FILLER_0_114_1003 ();
 sg13g2_fill_2 FILLER_0_114_1009 ();
 sg13g2_fill_8 FILLER_0_114_1016 ();
 sg13g2_fill_2 FILLER_0_114_1024 ();
 sg13g2_fill_1 FILLER_0_114_1026 ();
 sg13g2_fill_2 FILLER_0_114_1032 ();
 sg13g2_fill_8 FILLER_0_114_1039 ();
 sg13g2_fill_8 FILLER_0_114_1047 ();
 sg13g2_fill_8 FILLER_0_114_1055 ();
 sg13g2_fill_8 FILLER_0_114_1063 ();
 sg13g2_fill_1 FILLER_0_114_1071 ();
 sg13g2_fill_2 FILLER_0_114_1079 ();
 sg13g2_fill_8 FILLER_0_114_1086 ();
 sg13g2_fill_8 FILLER_0_114_1094 ();
 sg13g2_fill_2 FILLER_0_114_1107 ();
 sg13g2_fill_8 FILLER_0_114_1113 ();
 sg13g2_fill_8 FILLER_0_114_1121 ();
 sg13g2_fill_4 FILLER_0_114_1141 ();
 sg13g2_fill_2 FILLER_0_114_1145 ();
 sg13g2_fill_2 FILLER_0_114_1151 ();
 sg13g2_fill_8 FILLER_0_114_1157 ();
 sg13g2_fill_4 FILLER_0_114_1169 ();
 sg13g2_fill_2 FILLER_0_114_1173 ();
 sg13g2_fill_4 FILLER_0_114_1180 ();
 sg13g2_fill_2 FILLER_0_114_1184 ();
 sg13g2_fill_1 FILLER_0_114_1186 ();
 sg13g2_fill_2 FILLER_0_114_1197 ();
 sg13g2_fill_8 FILLER_0_114_1204 ();
 sg13g2_fill_8 FILLER_0_114_1212 ();
 sg13g2_fill_8 FILLER_0_114_1220 ();
 sg13g2_fill_8 FILLER_0_114_1228 ();
 sg13g2_fill_8 FILLER_0_114_1236 ();
 sg13g2_fill_1 FILLER_0_114_1244 ();
 sg13g2_fill_2 FILLER_0_114_1255 ();
 sg13g2_fill_1 FILLER_0_114_1257 ();
 sg13g2_fill_4 FILLER_0_114_1262 ();
 sg13g2_fill_1 FILLER_0_114_1266 ();
 sg13g2_fill_8 FILLER_0_114_1275 ();
 sg13g2_fill_2 FILLER_0_114_1286 ();
 sg13g2_fill_4 FILLER_0_114_1292 ();
 sg13g2_fill_1 FILLER_0_114_1296 ();
 sg13g2_fill_8 FILLER_0_115_0 ();
 sg13g2_fill_8 FILLER_0_115_8 ();
 sg13g2_fill_8 FILLER_0_115_16 ();
 sg13g2_fill_8 FILLER_0_115_24 ();
 sg13g2_fill_8 FILLER_0_115_32 ();
 sg13g2_fill_8 FILLER_0_115_40 ();
 sg13g2_fill_8 FILLER_0_115_48 ();
 sg13g2_fill_8 FILLER_0_115_56 ();
 sg13g2_fill_8 FILLER_0_115_64 ();
 sg13g2_fill_8 FILLER_0_115_72 ();
 sg13g2_fill_8 FILLER_0_115_80 ();
 sg13g2_fill_8 FILLER_0_115_88 ();
 sg13g2_fill_8 FILLER_0_115_96 ();
 sg13g2_fill_8 FILLER_0_115_104 ();
 sg13g2_fill_8 FILLER_0_115_112 ();
 sg13g2_fill_8 FILLER_0_115_120 ();
 sg13g2_fill_8 FILLER_0_115_128 ();
 sg13g2_fill_8 FILLER_0_115_136 ();
 sg13g2_fill_8 FILLER_0_115_144 ();
 sg13g2_fill_8 FILLER_0_115_152 ();
 sg13g2_fill_8 FILLER_0_115_160 ();
 sg13g2_fill_8 FILLER_0_115_168 ();
 sg13g2_fill_8 FILLER_0_115_176 ();
 sg13g2_fill_8 FILLER_0_115_184 ();
 sg13g2_fill_8 FILLER_0_115_192 ();
 sg13g2_fill_8 FILLER_0_115_200 ();
 sg13g2_fill_8 FILLER_0_115_208 ();
 sg13g2_fill_8 FILLER_0_115_216 ();
 sg13g2_fill_8 FILLER_0_115_224 ();
 sg13g2_fill_8 FILLER_0_115_232 ();
 sg13g2_fill_8 FILLER_0_115_240 ();
 sg13g2_fill_8 FILLER_0_115_248 ();
 sg13g2_fill_4 FILLER_0_115_256 ();
 sg13g2_fill_2 FILLER_0_115_266 ();
 sg13g2_fill_8 FILLER_0_115_273 ();
 sg13g2_fill_8 FILLER_0_115_281 ();
 sg13g2_fill_8 FILLER_0_115_289 ();
 sg13g2_fill_8 FILLER_0_115_297 ();
 sg13g2_fill_8 FILLER_0_115_305 ();
 sg13g2_fill_8 FILLER_0_115_313 ();
 sg13g2_fill_4 FILLER_0_115_321 ();
 sg13g2_fill_2 FILLER_0_115_325 ();
 sg13g2_fill_1 FILLER_0_115_327 ();
 sg13g2_fill_8 FILLER_0_115_354 ();
 sg13g2_fill_8 FILLER_0_115_362 ();
 sg13g2_fill_4 FILLER_0_115_370 ();
 sg13g2_fill_8 FILLER_0_115_379 ();
 sg13g2_fill_8 FILLER_0_115_387 ();
 sg13g2_fill_8 FILLER_0_115_395 ();
 sg13g2_fill_8 FILLER_0_115_403 ();
 sg13g2_fill_8 FILLER_0_115_411 ();
 sg13g2_fill_8 FILLER_0_115_419 ();
 sg13g2_fill_8 FILLER_0_115_427 ();
 sg13g2_fill_8 FILLER_0_115_435 ();
 sg13g2_fill_4 FILLER_0_115_443 ();
 sg13g2_fill_2 FILLER_0_115_451 ();
 sg13g2_fill_8 FILLER_0_115_458 ();
 sg13g2_fill_2 FILLER_0_115_471 ();
 sg13g2_fill_8 FILLER_0_115_481 ();
 sg13g2_fill_8 FILLER_0_115_489 ();
 sg13g2_fill_4 FILLER_0_115_497 ();
 sg13g2_fill_8 FILLER_0_115_506 ();
 sg13g2_fill_4 FILLER_0_115_514 ();
 sg13g2_fill_8 FILLER_0_115_523 ();
 sg13g2_fill_1 FILLER_0_115_531 ();
 sg13g2_fill_2 FILLER_0_115_537 ();
 sg13g2_fill_8 FILLER_0_115_543 ();
 sg13g2_fill_8 FILLER_0_115_551 ();
 sg13g2_fill_4 FILLER_0_115_559 ();
 sg13g2_fill_2 FILLER_0_115_563 ();
 sg13g2_fill_2 FILLER_0_115_571 ();
 sg13g2_fill_4 FILLER_0_115_579 ();
 sg13g2_fill_2 FILLER_0_115_583 ();
 sg13g2_fill_1 FILLER_0_115_585 ();
 sg13g2_fill_2 FILLER_0_115_590 ();
 sg13g2_fill_8 FILLER_0_115_618 ();
 sg13g2_fill_4 FILLER_0_115_626 ();
 sg13g2_fill_2 FILLER_0_115_630 ();
 sg13g2_fill_2 FILLER_0_115_636 ();
 sg13g2_fill_2 FILLER_0_115_642 ();
 sg13g2_fill_2 FILLER_0_115_649 ();
 sg13g2_fill_1 FILLER_0_115_651 ();
 sg13g2_fill_2 FILLER_0_115_657 ();
 sg13g2_fill_4 FILLER_0_115_664 ();
 sg13g2_fill_2 FILLER_0_115_673 ();
 sg13g2_fill_1 FILLER_0_115_675 ();
 sg13g2_fill_8 FILLER_0_115_681 ();
 sg13g2_fill_4 FILLER_0_115_689 ();
 sg13g2_fill_2 FILLER_0_115_693 ();
 sg13g2_fill_1 FILLER_0_115_695 ();
 sg13g2_fill_8 FILLER_0_115_702 ();
 sg13g2_fill_8 FILLER_0_115_710 ();
 sg13g2_fill_4 FILLER_0_115_718 ();
 sg13g2_fill_2 FILLER_0_115_722 ();
 sg13g2_fill_1 FILLER_0_115_724 ();
 sg13g2_fill_2 FILLER_0_115_730 ();
 sg13g2_fill_4 FILLER_0_115_736 ();
 sg13g2_fill_1 FILLER_0_115_740 ();
 sg13g2_fill_8 FILLER_0_115_751 ();
 sg13g2_fill_8 FILLER_0_115_759 ();
 sg13g2_fill_2 FILLER_0_115_767 ();
 sg13g2_fill_8 FILLER_0_115_774 ();
 sg13g2_fill_4 FILLER_0_115_782 ();
 sg13g2_fill_2 FILLER_0_115_786 ();
 sg13g2_fill_8 FILLER_0_115_814 ();
 sg13g2_fill_8 FILLER_0_115_822 ();
 sg13g2_fill_2 FILLER_0_115_834 ();
 sg13g2_fill_8 FILLER_0_115_841 ();
 sg13g2_fill_4 FILLER_0_115_870 ();
 sg13g2_fill_2 FILLER_0_115_874 ();
 sg13g2_fill_2 FILLER_0_115_881 ();
 sg13g2_fill_2 FILLER_0_115_888 ();
 sg13g2_fill_8 FILLER_0_115_895 ();
 sg13g2_fill_8 FILLER_0_115_908 ();
 sg13g2_fill_4 FILLER_0_115_916 ();
 sg13g2_fill_1 FILLER_0_115_920 ();
 sg13g2_fill_2 FILLER_0_115_925 ();
 sg13g2_fill_8 FILLER_0_115_932 ();
 sg13g2_fill_8 FILLER_0_115_940 ();
 sg13g2_fill_8 FILLER_0_115_948 ();
 sg13g2_fill_8 FILLER_0_115_956 ();
 sg13g2_fill_8 FILLER_0_115_964 ();
 sg13g2_fill_8 FILLER_0_115_972 ();
 sg13g2_fill_8 FILLER_0_115_980 ();
 sg13g2_fill_8 FILLER_0_115_988 ();
 sg13g2_fill_2 FILLER_0_115_996 ();
 sg13g2_fill_1 FILLER_0_115_998 ();
 sg13g2_fill_2 FILLER_0_115_1004 ();
 sg13g2_fill_8 FILLER_0_115_1011 ();
 sg13g2_fill_8 FILLER_0_115_1019 ();
 sg13g2_fill_2 FILLER_0_115_1027 ();
 sg13g2_fill_1 FILLER_0_115_1029 ();
 sg13g2_fill_2 FILLER_0_115_1038 ();
 sg13g2_fill_8 FILLER_0_115_1044 ();
 sg13g2_fill_8 FILLER_0_115_1052 ();
 sg13g2_fill_8 FILLER_0_115_1060 ();
 sg13g2_fill_8 FILLER_0_115_1068 ();
 sg13g2_fill_8 FILLER_0_115_1076 ();
 sg13g2_fill_8 FILLER_0_115_1084 ();
 sg13g2_fill_1 FILLER_0_115_1092 ();
 sg13g2_fill_2 FILLER_0_115_1101 ();
 sg13g2_fill_8 FILLER_0_115_1108 ();
 sg13g2_fill_2 FILLER_0_115_1124 ();
 sg13g2_fill_4 FILLER_0_115_1134 ();
 sg13g2_fill_8 FILLER_0_115_1146 ();
 sg13g2_fill_8 FILLER_0_115_1154 ();
 sg13g2_fill_1 FILLER_0_115_1162 ();
 sg13g2_fill_4 FILLER_0_115_1171 ();
 sg13g2_fill_2 FILLER_0_115_1175 ();
 sg13g2_fill_1 FILLER_0_115_1177 ();
 sg13g2_fill_4 FILLER_0_115_1182 ();
 sg13g2_fill_2 FILLER_0_115_1186 ();
 sg13g2_fill_8 FILLER_0_115_1193 ();
 sg13g2_fill_8 FILLER_0_115_1201 ();
 sg13g2_fill_8 FILLER_0_115_1209 ();
 sg13g2_fill_2 FILLER_0_115_1217 ();
 sg13g2_fill_1 FILLER_0_115_1219 ();
 sg13g2_fill_2 FILLER_0_115_1224 ();
 sg13g2_fill_4 FILLER_0_115_1230 ();
 sg13g2_fill_4 FILLER_0_115_1238 ();
 sg13g2_fill_1 FILLER_0_115_1242 ();
 sg13g2_fill_2 FILLER_0_115_1253 ();
 sg13g2_fill_2 FILLER_0_115_1281 ();
 sg13g2_fill_2 FILLER_0_115_1288 ();
 sg13g2_fill_1 FILLER_0_115_1290 ();
 sg13g2_fill_2 FILLER_0_115_1295 ();
 sg13g2_fill_8 FILLER_0_116_0 ();
 sg13g2_fill_8 FILLER_0_116_8 ();
 sg13g2_fill_8 FILLER_0_116_16 ();
 sg13g2_fill_8 FILLER_0_116_24 ();
 sg13g2_fill_8 FILLER_0_116_32 ();
 sg13g2_fill_8 FILLER_0_116_40 ();
 sg13g2_fill_8 FILLER_0_116_48 ();
 sg13g2_fill_8 FILLER_0_116_56 ();
 sg13g2_fill_8 FILLER_0_116_64 ();
 sg13g2_fill_8 FILLER_0_116_72 ();
 sg13g2_fill_8 FILLER_0_116_80 ();
 sg13g2_fill_8 FILLER_0_116_88 ();
 sg13g2_fill_8 FILLER_0_116_96 ();
 sg13g2_fill_8 FILLER_0_116_104 ();
 sg13g2_fill_8 FILLER_0_116_112 ();
 sg13g2_fill_8 FILLER_0_116_120 ();
 sg13g2_fill_8 FILLER_0_116_128 ();
 sg13g2_fill_8 FILLER_0_116_136 ();
 sg13g2_fill_8 FILLER_0_116_144 ();
 sg13g2_fill_8 FILLER_0_116_152 ();
 sg13g2_fill_8 FILLER_0_116_160 ();
 sg13g2_fill_8 FILLER_0_116_168 ();
 sg13g2_fill_8 FILLER_0_116_176 ();
 sg13g2_fill_8 FILLER_0_116_184 ();
 sg13g2_fill_8 FILLER_0_116_192 ();
 sg13g2_fill_8 FILLER_0_116_200 ();
 sg13g2_fill_4 FILLER_0_116_208 ();
 sg13g2_fill_2 FILLER_0_116_212 ();
 sg13g2_fill_8 FILLER_0_116_219 ();
 sg13g2_fill_1 FILLER_0_116_227 ();
 sg13g2_fill_8 FILLER_0_116_232 ();
 sg13g2_fill_4 FILLER_0_116_240 ();
 sg13g2_fill_4 FILLER_0_116_249 ();
 sg13g2_fill_2 FILLER_0_116_253 ();
 sg13g2_fill_1 FILLER_0_116_255 ();
 sg13g2_fill_4 FILLER_0_116_262 ();
 sg13g2_fill_2 FILLER_0_116_266 ();
 sg13g2_fill_1 FILLER_0_116_268 ();
 sg13g2_fill_2 FILLER_0_116_274 ();
 sg13g2_fill_2 FILLER_0_116_281 ();
 sg13g2_fill_8 FILLER_0_116_289 ();
 sg13g2_fill_2 FILLER_0_116_297 ();
 sg13g2_fill_2 FILLER_0_116_304 ();
 sg13g2_fill_2 FILLER_0_116_310 ();
 sg13g2_fill_1 FILLER_0_116_312 ();
 sg13g2_fill_8 FILLER_0_116_317 ();
 sg13g2_fill_8 FILLER_0_116_325 ();
 sg13g2_fill_8 FILLER_0_116_337 ();
 sg13g2_fill_4 FILLER_0_116_345 ();
 sg13g2_fill_1 FILLER_0_116_349 ();
 sg13g2_fill_8 FILLER_0_116_355 ();
 sg13g2_fill_8 FILLER_0_116_363 ();
 sg13g2_fill_8 FILLER_0_116_371 ();
 sg13g2_fill_8 FILLER_0_116_379 ();
 sg13g2_fill_8 FILLER_0_116_387 ();
 sg13g2_fill_8 FILLER_0_116_395 ();
 sg13g2_fill_8 FILLER_0_116_403 ();
 sg13g2_fill_8 FILLER_0_116_411 ();
 sg13g2_fill_8 FILLER_0_116_419 ();
 sg13g2_fill_8 FILLER_0_116_427 ();
 sg13g2_fill_8 FILLER_0_116_435 ();
 sg13g2_fill_4 FILLER_0_116_443 ();
 sg13g2_fill_2 FILLER_0_116_455 ();
 sg13g2_fill_4 FILLER_0_116_461 ();
 sg13g2_fill_2 FILLER_0_116_465 ();
 sg13g2_fill_1 FILLER_0_116_467 ();
 sg13g2_fill_2 FILLER_0_116_473 ();
 sg13g2_fill_8 FILLER_0_116_479 ();
 sg13g2_fill_8 FILLER_0_116_487 ();
 sg13g2_fill_4 FILLER_0_116_495 ();
 sg13g2_fill_2 FILLER_0_116_499 ();
 sg13g2_fill_8 FILLER_0_116_506 ();
 sg13g2_fill_1 FILLER_0_116_514 ();
 sg13g2_fill_8 FILLER_0_116_541 ();
 sg13g2_fill_8 FILLER_0_116_549 ();
 sg13g2_fill_8 FILLER_0_116_557 ();
 sg13g2_fill_8 FILLER_0_116_565 ();
 sg13g2_fill_8 FILLER_0_116_573 ();
 sg13g2_fill_2 FILLER_0_116_581 ();
 sg13g2_fill_1 FILLER_0_116_583 ();
 sg13g2_fill_8 FILLER_0_116_589 ();
 sg13g2_fill_8 FILLER_0_116_602 ();
 sg13g2_fill_2 FILLER_0_116_615 ();
 sg13g2_fill_4 FILLER_0_116_622 ();
 sg13g2_fill_1 FILLER_0_116_626 ();
 sg13g2_fill_2 FILLER_0_116_632 ();
 sg13g2_fill_2 FILLER_0_116_639 ();
 sg13g2_fill_2 FILLER_0_116_667 ();
 sg13g2_fill_2 FILLER_0_116_674 ();
 sg13g2_fill_8 FILLER_0_116_681 ();
 sg13g2_fill_4 FILLER_0_116_689 ();
 sg13g2_fill_2 FILLER_0_116_693 ();
 sg13g2_fill_1 FILLER_0_116_695 ();
 sg13g2_fill_4 FILLER_0_116_701 ();
 sg13g2_fill_8 FILLER_0_116_709 ();
 sg13g2_fill_8 FILLER_0_116_717 ();
 sg13g2_fill_1 FILLER_0_116_725 ();
 sg13g2_fill_8 FILLER_0_116_730 ();
 sg13g2_fill_4 FILLER_0_116_738 ();
 sg13g2_fill_2 FILLER_0_116_742 ();
 sg13g2_fill_8 FILLER_0_116_749 ();
 sg13g2_fill_8 FILLER_0_116_757 ();
 sg13g2_fill_4 FILLER_0_116_765 ();
 sg13g2_fill_8 FILLER_0_116_774 ();
 sg13g2_fill_8 FILLER_0_116_782 ();
 sg13g2_fill_2 FILLER_0_116_790 ();
 sg13g2_fill_2 FILLER_0_116_797 ();
 sg13g2_fill_2 FILLER_0_116_803 ();
 sg13g2_fill_2 FILLER_0_116_810 ();
 sg13g2_fill_8 FILLER_0_116_817 ();
 sg13g2_fill_1 FILLER_0_116_825 ();
 sg13g2_fill_8 FILLER_0_116_830 ();
 sg13g2_fill_8 FILLER_0_116_838 ();
 sg13g2_fill_4 FILLER_0_116_846 ();
 sg13g2_fill_1 FILLER_0_116_850 ();
 sg13g2_fill_2 FILLER_0_116_855 ();
 sg13g2_fill_2 FILLER_0_116_862 ();
 sg13g2_fill_1 FILLER_0_116_864 ();
 sg13g2_fill_4 FILLER_0_116_869 ();
 sg13g2_fill_2 FILLER_0_116_877 ();
 sg13g2_fill_1 FILLER_0_116_879 ();
 sg13g2_fill_8 FILLER_0_116_885 ();
 sg13g2_fill_8 FILLER_0_116_893 ();
 sg13g2_fill_8 FILLER_0_116_901 ();
 sg13g2_fill_8 FILLER_0_116_909 ();
 sg13g2_fill_8 FILLER_0_116_917 ();
 sg13g2_fill_4 FILLER_0_116_925 ();
 sg13g2_fill_8 FILLER_0_116_933 ();
 sg13g2_fill_8 FILLER_0_116_941 ();
 sg13g2_fill_4 FILLER_0_116_949 ();
 sg13g2_fill_2 FILLER_0_116_953 ();
 sg13g2_fill_1 FILLER_0_116_955 ();
 sg13g2_fill_8 FILLER_0_116_961 ();
 sg13g2_fill_8 FILLER_0_116_969 ();
 sg13g2_fill_8 FILLER_0_116_977 ();
 sg13g2_fill_8 FILLER_0_116_985 ();
 sg13g2_fill_1 FILLER_0_116_993 ();
 sg13g2_fill_2 FILLER_0_116_1002 ();
 sg13g2_fill_2 FILLER_0_116_1008 ();
 sg13g2_fill_8 FILLER_0_116_1015 ();
 sg13g2_fill_8 FILLER_0_116_1023 ();
 sg13g2_fill_2 FILLER_0_116_1031 ();
 sg13g2_fill_2 FILLER_0_116_1037 ();
 sg13g2_fill_4 FILLER_0_116_1043 ();
 sg13g2_fill_8 FILLER_0_116_1052 ();
 sg13g2_fill_8 FILLER_0_116_1060 ();
 sg13g2_fill_4 FILLER_0_116_1068 ();
 sg13g2_fill_1 FILLER_0_116_1072 ();
 sg13g2_fill_8 FILLER_0_116_1080 ();
 sg13g2_fill_8 FILLER_0_116_1088 ();
 sg13g2_fill_1 FILLER_0_116_1096 ();
 sg13g2_fill_2 FILLER_0_116_1101 ();
 sg13g2_fill_2 FILLER_0_116_1108 ();
 sg13g2_fill_2 FILLER_0_116_1117 ();
 sg13g2_fill_2 FILLER_0_116_1124 ();
 sg13g2_fill_2 FILLER_0_116_1130 ();
 sg13g2_fill_1 FILLER_0_116_1132 ();
 sg13g2_fill_8 FILLER_0_116_1138 ();
 sg13g2_fill_4 FILLER_0_116_1146 ();
 sg13g2_fill_2 FILLER_0_116_1150 ();
 sg13g2_fill_8 FILLER_0_116_1161 ();
 sg13g2_fill_8 FILLER_0_116_1169 ();
 sg13g2_fill_4 FILLER_0_116_1177 ();
 sg13g2_fill_2 FILLER_0_116_1181 ();
 sg13g2_fill_8 FILLER_0_116_1187 ();
 sg13g2_fill_8 FILLER_0_116_1195 ();
 sg13g2_fill_8 FILLER_0_116_1203 ();
 sg13g2_fill_2 FILLER_0_116_1211 ();
 sg13g2_fill_2 FILLER_0_116_1217 ();
 sg13g2_fill_2 FILLER_0_116_1224 ();
 sg13g2_fill_2 FILLER_0_116_1231 ();
 sg13g2_fill_8 FILLER_0_116_1238 ();
 sg13g2_fill_8 FILLER_0_116_1246 ();
 sg13g2_fill_2 FILLER_0_116_1254 ();
 sg13g2_fill_4 FILLER_0_116_1260 ();
 sg13g2_fill_8 FILLER_0_116_1268 ();
 sg13g2_fill_1 FILLER_0_116_1276 ();
 sg13g2_fill_2 FILLER_0_116_1281 ();
 sg13g2_fill_4 FILLER_0_116_1287 ();
 sg13g2_fill_1 FILLER_0_116_1291 ();
 sg13g2_fill_1 FILLER_0_116_1296 ();
 sg13g2_fill_8 FILLER_0_117_0 ();
 sg13g2_fill_8 FILLER_0_117_8 ();
 sg13g2_fill_8 FILLER_0_117_16 ();
 sg13g2_fill_8 FILLER_0_117_24 ();
 sg13g2_fill_8 FILLER_0_117_32 ();
 sg13g2_fill_8 FILLER_0_117_40 ();
 sg13g2_fill_8 FILLER_0_117_48 ();
 sg13g2_fill_8 FILLER_0_117_56 ();
 sg13g2_fill_8 FILLER_0_117_64 ();
 sg13g2_fill_8 FILLER_0_117_72 ();
 sg13g2_fill_8 FILLER_0_117_80 ();
 sg13g2_fill_8 FILLER_0_117_88 ();
 sg13g2_fill_8 FILLER_0_117_96 ();
 sg13g2_fill_8 FILLER_0_117_104 ();
 sg13g2_fill_8 FILLER_0_117_112 ();
 sg13g2_fill_8 FILLER_0_117_120 ();
 sg13g2_fill_8 FILLER_0_117_128 ();
 sg13g2_fill_8 FILLER_0_117_136 ();
 sg13g2_fill_8 FILLER_0_117_144 ();
 sg13g2_fill_8 FILLER_0_117_152 ();
 sg13g2_fill_8 FILLER_0_117_160 ();
 sg13g2_fill_8 FILLER_0_117_168 ();
 sg13g2_fill_8 FILLER_0_117_176 ();
 sg13g2_fill_8 FILLER_0_117_184 ();
 sg13g2_fill_8 FILLER_0_117_192 ();
 sg13g2_fill_8 FILLER_0_117_200 ();
 sg13g2_fill_2 FILLER_0_117_208 ();
 sg13g2_fill_1 FILLER_0_117_210 ();
 sg13g2_fill_8 FILLER_0_117_237 ();
 sg13g2_fill_2 FILLER_0_117_245 ();
 sg13g2_fill_1 FILLER_0_117_247 ();
 sg13g2_fill_4 FILLER_0_117_274 ();
 sg13g2_fill_2 FILLER_0_117_283 ();
 sg13g2_fill_1 FILLER_0_117_285 ();
 sg13g2_fill_4 FILLER_0_117_294 ();
 sg13g2_fill_8 FILLER_0_117_324 ();
 sg13g2_fill_8 FILLER_0_117_332 ();
 sg13g2_fill_8 FILLER_0_117_340 ();
 sg13g2_fill_2 FILLER_0_117_348 ();
 sg13g2_fill_8 FILLER_0_117_376 ();
 sg13g2_fill_8 FILLER_0_117_384 ();
 sg13g2_fill_2 FILLER_0_117_392 ();
 sg13g2_fill_1 FILLER_0_117_394 ();
 sg13g2_fill_2 FILLER_0_117_400 ();
 sg13g2_fill_4 FILLER_0_117_406 ();
 sg13g2_fill_2 FILLER_0_117_410 ();
 sg13g2_fill_2 FILLER_0_117_416 ();
 sg13g2_fill_1 FILLER_0_117_418 ();
 sg13g2_fill_8 FILLER_0_117_427 ();
 sg13g2_fill_8 FILLER_0_117_435 ();
 sg13g2_fill_8 FILLER_0_117_443 ();
 sg13g2_fill_2 FILLER_0_117_451 ();
 sg13g2_fill_8 FILLER_0_117_458 ();
 sg13g2_fill_4 FILLER_0_117_466 ();
 sg13g2_fill_2 FILLER_0_117_470 ();
 sg13g2_fill_1 FILLER_0_117_472 ();
 sg13g2_fill_2 FILLER_0_117_499 ();
 sg13g2_fill_8 FILLER_0_117_506 ();
 sg13g2_fill_8 FILLER_0_117_514 ();
 sg13g2_fill_8 FILLER_0_117_522 ();
 sg13g2_fill_2 FILLER_0_117_530 ();
 sg13g2_fill_8 FILLER_0_117_537 ();
 sg13g2_fill_1 FILLER_0_117_545 ();
 sg13g2_fill_2 FILLER_0_117_550 ();
 sg13g2_fill_8 FILLER_0_117_562 ();
 sg13g2_fill_8 FILLER_0_117_570 ();
 sg13g2_fill_8 FILLER_0_117_578 ();
 sg13g2_fill_8 FILLER_0_117_586 ();
 sg13g2_fill_8 FILLER_0_117_594 ();
 sg13g2_fill_8 FILLER_0_117_602 ();
 sg13g2_fill_8 FILLER_0_117_610 ();
 sg13g2_fill_8 FILLER_0_117_618 ();
 sg13g2_fill_8 FILLER_0_117_626 ();
 sg13g2_fill_8 FILLER_0_117_634 ();
 sg13g2_fill_8 FILLER_0_117_642 ();
 sg13g2_fill_2 FILLER_0_117_655 ();
 sg13g2_fill_8 FILLER_0_117_678 ();
 sg13g2_fill_4 FILLER_0_117_686 ();
 sg13g2_fill_8 FILLER_0_117_716 ();
 sg13g2_fill_4 FILLER_0_117_724 ();
 sg13g2_fill_1 FILLER_0_117_728 ();
 sg13g2_fill_8 FILLER_0_117_734 ();
 sg13g2_fill_2 FILLER_0_117_742 ();
 sg13g2_fill_1 FILLER_0_117_744 ();
 sg13g2_fill_8 FILLER_0_117_753 ();
 sg13g2_fill_8 FILLER_0_117_761 ();
 sg13g2_fill_8 FILLER_0_117_769 ();
 sg13g2_fill_2 FILLER_0_117_782 ();
 sg13g2_fill_4 FILLER_0_117_788 ();
 sg13g2_fill_2 FILLER_0_117_792 ();
 sg13g2_fill_2 FILLER_0_117_804 ();
 sg13g2_fill_4 FILLER_0_117_811 ();
 sg13g2_fill_2 FILLER_0_117_815 ();
 sg13g2_fill_1 FILLER_0_117_817 ();
 sg13g2_fill_2 FILLER_0_117_822 ();
 sg13g2_fill_2 FILLER_0_117_828 ();
 sg13g2_fill_2 FILLER_0_117_836 ();
 sg13g2_fill_4 FILLER_0_117_846 ();
 sg13g2_fill_1 FILLER_0_117_850 ();
 sg13g2_fill_2 FILLER_0_117_877 ();
 sg13g2_fill_8 FILLER_0_117_884 ();
 sg13g2_fill_8 FILLER_0_117_892 ();
 sg13g2_fill_4 FILLER_0_117_900 ();
 sg13g2_fill_2 FILLER_0_117_904 ();
 sg13g2_fill_1 FILLER_0_117_906 ();
 sg13g2_fill_2 FILLER_0_117_912 ();
 sg13g2_fill_4 FILLER_0_117_919 ();
 sg13g2_fill_1 FILLER_0_117_923 ();
 sg13g2_fill_2 FILLER_0_117_928 ();
 sg13g2_fill_2 FILLER_0_117_936 ();
 sg13g2_fill_2 FILLER_0_117_943 ();
 sg13g2_fill_2 FILLER_0_117_950 ();
 sg13g2_fill_2 FILLER_0_117_956 ();
 sg13g2_fill_4 FILLER_0_117_963 ();
 sg13g2_fill_8 FILLER_0_117_973 ();
 sg13g2_fill_4 FILLER_0_117_981 ();
 sg13g2_fill_2 FILLER_0_117_985 ();
 sg13g2_fill_1 FILLER_0_117_987 ();
 sg13g2_fill_8 FILLER_0_117_992 ();
 sg13g2_fill_8 FILLER_0_117_1000 ();
 sg13g2_fill_8 FILLER_0_117_1008 ();
 sg13g2_fill_2 FILLER_0_117_1021 ();
 sg13g2_fill_4 FILLER_0_117_1027 ();
 sg13g2_fill_2 FILLER_0_117_1037 ();
 sg13g2_fill_8 FILLER_0_117_1043 ();
 sg13g2_fill_4 FILLER_0_117_1051 ();
 sg13g2_fill_1 FILLER_0_117_1055 ();
 sg13g2_fill_4 FILLER_0_117_1062 ();
 sg13g2_fill_2 FILLER_0_117_1066 ();
 sg13g2_fill_1 FILLER_0_117_1068 ();
 sg13g2_fill_2 FILLER_0_117_1075 ();
 sg13g2_fill_8 FILLER_0_117_1085 ();
 sg13g2_fill_8 FILLER_0_117_1093 ();
 sg13g2_fill_8 FILLER_0_117_1101 ();
 sg13g2_fill_2 FILLER_0_117_1109 ();
 sg13g2_fill_2 FILLER_0_117_1114 ();
 sg13g2_fill_2 FILLER_0_117_1121 ();
 sg13g2_fill_8 FILLER_0_117_1128 ();
 sg13g2_fill_2 FILLER_0_117_1140 ();
 sg13g2_fill_4 FILLER_0_117_1146 ();
 sg13g2_fill_2 FILLER_0_117_1150 ();
 sg13g2_fill_8 FILLER_0_117_1158 ();
 sg13g2_fill_2 FILLER_0_117_1166 ();
 sg13g2_fill_1 FILLER_0_117_1168 ();
 sg13g2_fill_2 FILLER_0_117_1175 ();
 sg13g2_fill_2 FILLER_0_117_1182 ();
 sg13g2_fill_2 FILLER_0_117_1190 ();
 sg13g2_fill_2 FILLER_0_117_1197 ();
 sg13g2_fill_2 FILLER_0_117_1203 ();
 sg13g2_fill_2 FILLER_0_117_1210 ();
 sg13g2_fill_1 FILLER_0_117_1212 ();
 sg13g2_fill_2 FILLER_0_117_1218 ();
 sg13g2_fill_2 FILLER_0_117_1226 ();
 sg13g2_fill_1 FILLER_0_117_1228 ();
 sg13g2_fill_2 FILLER_0_117_1233 ();
 sg13g2_fill_8 FILLER_0_117_1239 ();
 sg13g2_fill_1 FILLER_0_117_1247 ();
 sg13g2_fill_2 FILLER_0_117_1252 ();
 sg13g2_fill_2 FILLER_0_117_1259 ();
 sg13g2_fill_4 FILLER_0_117_1265 ();
 sg13g2_fill_2 FILLER_0_117_1269 ();
 sg13g2_fill_1 FILLER_0_117_1271 ();
 sg13g2_fill_2 FILLER_0_117_1276 ();
 sg13g2_fill_2 FILLER_0_117_1282 ();
 sg13g2_fill_2 FILLER_0_117_1288 ();
 sg13g2_fill_2 FILLER_0_117_1294 ();
 sg13g2_fill_1 FILLER_0_117_1296 ();
 sg13g2_fill_8 FILLER_0_118_0 ();
 sg13g2_fill_8 FILLER_0_118_8 ();
 sg13g2_fill_8 FILLER_0_118_16 ();
 sg13g2_fill_8 FILLER_0_118_24 ();
 sg13g2_fill_8 FILLER_0_118_32 ();
 sg13g2_fill_8 FILLER_0_118_40 ();
 sg13g2_fill_8 FILLER_0_118_48 ();
 sg13g2_fill_8 FILLER_0_118_56 ();
 sg13g2_fill_8 FILLER_0_118_64 ();
 sg13g2_fill_8 FILLER_0_118_72 ();
 sg13g2_fill_8 FILLER_0_118_80 ();
 sg13g2_fill_8 FILLER_0_118_88 ();
 sg13g2_fill_8 FILLER_0_118_96 ();
 sg13g2_fill_8 FILLER_0_118_104 ();
 sg13g2_fill_8 FILLER_0_118_112 ();
 sg13g2_fill_8 FILLER_0_118_120 ();
 sg13g2_fill_8 FILLER_0_118_128 ();
 sg13g2_fill_8 FILLER_0_118_136 ();
 sg13g2_fill_8 FILLER_0_118_144 ();
 sg13g2_fill_8 FILLER_0_118_152 ();
 sg13g2_fill_8 FILLER_0_118_160 ();
 sg13g2_fill_8 FILLER_0_118_168 ();
 sg13g2_fill_8 FILLER_0_118_176 ();
 sg13g2_fill_8 FILLER_0_118_184 ();
 sg13g2_fill_8 FILLER_0_118_192 ();
 sg13g2_fill_8 FILLER_0_118_200 ();
 sg13g2_fill_8 FILLER_0_118_208 ();
 sg13g2_fill_4 FILLER_0_118_216 ();
 sg13g2_fill_1 FILLER_0_118_220 ();
 sg13g2_fill_2 FILLER_0_118_247 ();
 sg13g2_fill_2 FILLER_0_118_255 ();
 sg13g2_fill_2 FILLER_0_118_263 ();
 sg13g2_fill_8 FILLER_0_118_269 ();
 sg13g2_fill_8 FILLER_0_118_277 ();
 sg13g2_fill_1 FILLER_0_118_285 ();
 sg13g2_fill_2 FILLER_0_118_292 ();
 sg13g2_fill_4 FILLER_0_118_299 ();
 sg13g2_fill_1 FILLER_0_118_303 ();
 sg13g2_fill_8 FILLER_0_118_309 ();
 sg13g2_fill_4 FILLER_0_118_317 ();
 sg13g2_fill_2 FILLER_0_118_326 ();
 sg13g2_fill_2 FILLER_0_118_333 ();
 sg13g2_fill_4 FILLER_0_118_340 ();
 sg13g2_fill_4 FILLER_0_118_350 ();
 sg13g2_fill_2 FILLER_0_118_354 ();
 sg13g2_fill_1 FILLER_0_118_356 ();
 sg13g2_fill_2 FILLER_0_118_362 ();
 sg13g2_fill_4 FILLER_0_118_390 ();
 sg13g2_fill_2 FILLER_0_118_399 ();
 sg13g2_fill_8 FILLER_0_118_427 ();
 sg13g2_fill_4 FILLER_0_118_435 ();
 sg13g2_fill_1 FILLER_0_118_439 ();
 sg13g2_fill_4 FILLER_0_118_466 ();
 sg13g2_fill_2 FILLER_0_118_470 ();
 sg13g2_fill_1 FILLER_0_118_472 ();
 sg13g2_fill_8 FILLER_0_118_478 ();
 sg13g2_fill_1 FILLER_0_118_486 ();
 sg13g2_fill_2 FILLER_0_118_492 ();
 sg13g2_fill_1 FILLER_0_118_494 ();
 sg13g2_fill_2 FILLER_0_118_500 ();
 sg13g2_fill_8 FILLER_0_118_510 ();
 sg13g2_fill_1 FILLER_0_118_518 ();
 sg13g2_fill_8 FILLER_0_118_524 ();
 sg13g2_fill_1 FILLER_0_118_532 ();
 sg13g2_fill_2 FILLER_0_118_559 ();
 sg13g2_fill_8 FILLER_0_118_566 ();
 sg13g2_fill_8 FILLER_0_118_579 ();
 sg13g2_fill_4 FILLER_0_118_587 ();
 sg13g2_fill_2 FILLER_0_118_596 ();
 sg13g2_fill_8 FILLER_0_118_602 ();
 sg13g2_fill_8 FILLER_0_118_610 ();
 sg13g2_fill_8 FILLER_0_118_618 ();
 sg13g2_fill_8 FILLER_0_118_626 ();
 sg13g2_fill_8 FILLER_0_118_634 ();
 sg13g2_fill_4 FILLER_0_118_642 ();
 sg13g2_fill_2 FILLER_0_118_646 ();
 sg13g2_fill_4 FILLER_0_118_674 ();
 sg13g2_fill_2 FILLER_0_118_683 ();
 sg13g2_fill_8 FILLER_0_118_693 ();
 sg13g2_fill_1 FILLER_0_118_701 ();
 sg13g2_fill_8 FILLER_0_118_710 ();
 sg13g2_fill_8 FILLER_0_118_728 ();
 sg13g2_fill_8 FILLER_0_118_736 ();
 sg13g2_fill_8 FILLER_0_118_744 ();
 sg13g2_fill_4 FILLER_0_118_752 ();
 sg13g2_fill_2 FILLER_0_118_756 ();
 sg13g2_fill_2 FILLER_0_118_784 ();
 sg13g2_fill_4 FILLER_0_118_796 ();
 sg13g2_fill_8 FILLER_0_118_805 ();
 sg13g2_fill_4 FILLER_0_118_813 ();
 sg13g2_fill_4 FILLER_0_118_825 ();
 sg13g2_fill_2 FILLER_0_118_829 ();
 sg13g2_fill_1 FILLER_0_118_831 ();
 sg13g2_fill_8 FILLER_0_118_858 ();
 sg13g2_fill_4 FILLER_0_118_866 ();
 sg13g2_fill_1 FILLER_0_118_870 ();
 sg13g2_fill_2 FILLER_0_118_881 ();
 sg13g2_fill_2 FILLER_0_118_887 ();
 sg13g2_fill_1 FILLER_0_118_889 ();
 sg13g2_fill_8 FILLER_0_118_894 ();
 sg13g2_fill_8 FILLER_0_118_902 ();
 sg13g2_fill_4 FILLER_0_118_910 ();
 sg13g2_fill_2 FILLER_0_118_914 ();
 sg13g2_fill_1 FILLER_0_118_916 ();
 sg13g2_fill_4 FILLER_0_118_922 ();
 sg13g2_fill_2 FILLER_0_118_926 ();
 sg13g2_fill_1 FILLER_0_118_928 ();
 sg13g2_fill_2 FILLER_0_118_936 ();
 sg13g2_fill_4 FILLER_0_118_946 ();
 sg13g2_fill_2 FILLER_0_118_950 ();
 sg13g2_fill_1 FILLER_0_118_952 ();
 sg13g2_fill_2 FILLER_0_118_958 ();
 sg13g2_fill_1 FILLER_0_118_960 ();
 sg13g2_fill_2 FILLER_0_118_968 ();
 sg13g2_fill_4 FILLER_0_118_975 ();
 sg13g2_fill_2 FILLER_0_118_984 ();
 sg13g2_fill_4 FILLER_0_118_992 ();
 sg13g2_fill_2 FILLER_0_118_996 ();
 sg13g2_fill_4 FILLER_0_118_1003 ();
 sg13g2_fill_1 FILLER_0_118_1007 ();
 sg13g2_fill_2 FILLER_0_118_1012 ();
 sg13g2_fill_2 FILLER_0_118_1020 ();
 sg13g2_fill_2 FILLER_0_118_1030 ();
 sg13g2_fill_2 FILLER_0_118_1037 ();
 sg13g2_fill_1 FILLER_0_118_1039 ();
 sg13g2_fill_2 FILLER_0_118_1046 ();
 sg13g2_fill_2 FILLER_0_118_1054 ();
 sg13g2_fill_2 FILLER_0_118_1062 ();
 sg13g2_fill_1 FILLER_0_118_1064 ();
 sg13g2_fill_8 FILLER_0_118_1071 ();
 sg13g2_fill_8 FILLER_0_118_1079 ();
 sg13g2_fill_8 FILLER_0_118_1087 ();
 sg13g2_fill_8 FILLER_0_118_1103 ();
 sg13g2_fill_1 FILLER_0_118_1111 ();
 sg13g2_fill_2 FILLER_0_118_1116 ();
 sg13g2_fill_2 FILLER_0_118_1123 ();
 sg13g2_fill_1 FILLER_0_118_1125 ();
 sg13g2_fill_4 FILLER_0_118_1134 ();
 sg13g2_fill_1 FILLER_0_118_1138 ();
 sg13g2_fill_8 FILLER_0_118_1144 ();
 sg13g2_fill_8 FILLER_0_118_1152 ();
 sg13g2_fill_4 FILLER_0_118_1160 ();
 sg13g2_fill_2 FILLER_0_118_1169 ();
 sg13g2_fill_2 FILLER_0_118_1179 ();
 sg13g2_fill_2 FILLER_0_118_1186 ();
 sg13g2_fill_4 FILLER_0_118_1193 ();
 sg13g2_fill_2 FILLER_0_118_1197 ();
 sg13g2_fill_1 FILLER_0_118_1199 ();
 sg13g2_fill_4 FILLER_0_118_1205 ();
 sg13g2_fill_1 FILLER_0_118_1209 ();
 sg13g2_fill_2 FILLER_0_118_1215 ();
 sg13g2_fill_2 FILLER_0_118_1222 ();
 sg13g2_fill_2 FILLER_0_118_1228 ();
 sg13g2_fill_2 FILLER_0_118_1235 ();
 sg13g2_fill_8 FILLER_0_118_1243 ();
 sg13g2_fill_4 FILLER_0_118_1251 ();
 sg13g2_fill_2 FILLER_0_118_1255 ();
 sg13g2_fill_8 FILLER_0_118_1261 ();
 sg13g2_fill_2 FILLER_0_118_1269 ();
 sg13g2_fill_4 FILLER_0_118_1275 ();
 sg13g2_fill_8 FILLER_0_118_1283 ();
 sg13g2_fill_4 FILLER_0_118_1291 ();
 sg13g2_fill_2 FILLER_0_118_1295 ();
 sg13g2_fill_8 FILLER_0_119_0 ();
 sg13g2_fill_8 FILLER_0_119_8 ();
 sg13g2_fill_4 FILLER_0_119_16 ();
 sg13g2_fill_8 FILLER_0_119_24 ();
 sg13g2_fill_8 FILLER_0_119_32 ();
 sg13g2_fill_8 FILLER_0_119_40 ();
 sg13g2_fill_8 FILLER_0_119_48 ();
 sg13g2_fill_8 FILLER_0_119_56 ();
 sg13g2_fill_8 FILLER_0_119_64 ();
 sg13g2_fill_8 FILLER_0_119_72 ();
 sg13g2_fill_8 FILLER_0_119_80 ();
 sg13g2_fill_8 FILLER_0_119_88 ();
 sg13g2_fill_8 FILLER_0_119_96 ();
 sg13g2_fill_8 FILLER_0_119_104 ();
 sg13g2_fill_8 FILLER_0_119_112 ();
 sg13g2_fill_8 FILLER_0_119_120 ();
 sg13g2_fill_8 FILLER_0_119_128 ();
 sg13g2_fill_8 FILLER_0_119_136 ();
 sg13g2_fill_8 FILLER_0_119_144 ();
 sg13g2_fill_8 FILLER_0_119_152 ();
 sg13g2_fill_8 FILLER_0_119_160 ();
 sg13g2_fill_8 FILLER_0_119_168 ();
 sg13g2_fill_8 FILLER_0_119_176 ();
 sg13g2_fill_8 FILLER_0_119_184 ();
 sg13g2_fill_8 FILLER_0_119_192 ();
 sg13g2_fill_8 FILLER_0_119_200 ();
 sg13g2_fill_8 FILLER_0_119_208 ();
 sg13g2_fill_4 FILLER_0_119_216 ();
 sg13g2_fill_2 FILLER_0_119_220 ();
 sg13g2_fill_1 FILLER_0_119_222 ();
 sg13g2_fill_8 FILLER_0_119_228 ();
 sg13g2_fill_4 FILLER_0_119_240 ();
 sg13g2_fill_2 FILLER_0_119_244 ();
 sg13g2_fill_1 FILLER_0_119_246 ();
 sg13g2_fill_8 FILLER_0_119_252 ();
 sg13g2_fill_8 FILLER_0_119_260 ();
 sg13g2_fill_8 FILLER_0_119_268 ();
 sg13g2_fill_8 FILLER_0_119_276 ();
 sg13g2_fill_8 FILLER_0_119_284 ();
 sg13g2_fill_8 FILLER_0_119_292 ();
 sg13g2_fill_8 FILLER_0_119_300 ();
 sg13g2_fill_2 FILLER_0_119_308 ();
 sg13g2_fill_2 FILLER_0_119_318 ();
 sg13g2_fill_2 FILLER_0_119_325 ();
 sg13g2_fill_8 FILLER_0_119_334 ();
 sg13g2_fill_2 FILLER_0_119_350 ();
 sg13g2_fill_2 FILLER_0_119_360 ();
 sg13g2_fill_2 FILLER_0_119_366 ();
 sg13g2_fill_2 FILLER_0_119_389 ();
 sg13g2_fill_2 FILLER_0_119_396 ();
 sg13g2_fill_4 FILLER_0_119_403 ();
 sg13g2_fill_2 FILLER_0_119_415 ();
 sg13g2_fill_4 FILLER_0_119_421 ();
 sg13g2_fill_1 FILLER_0_119_425 ();
 sg13g2_fill_2 FILLER_0_119_431 ();
 sg13g2_fill_4 FILLER_0_119_439 ();
 sg13g2_fill_2 FILLER_0_119_443 ();
 sg13g2_fill_1 FILLER_0_119_445 ();
 sg13g2_fill_2 FILLER_0_119_451 ();
 sg13g2_fill_1 FILLER_0_119_453 ();
 sg13g2_fill_2 FILLER_0_119_458 ();
 sg13g2_fill_4 FILLER_0_119_464 ();
 sg13g2_fill_8 FILLER_0_119_478 ();
 sg13g2_fill_8 FILLER_0_119_486 ();
 sg13g2_fill_4 FILLER_0_119_494 ();
 sg13g2_fill_2 FILLER_0_119_498 ();
 sg13g2_fill_1 FILLER_0_119_500 ();
 sg13g2_fill_8 FILLER_0_119_505 ();
 sg13g2_fill_8 FILLER_0_119_513 ();
 sg13g2_fill_4 FILLER_0_119_521 ();
 sg13g2_fill_2 FILLER_0_119_525 ();
 sg13g2_fill_1 FILLER_0_119_527 ();
 sg13g2_fill_8 FILLER_0_119_549 ();
 sg13g2_fill_1 FILLER_0_119_557 ();
 sg13g2_fill_2 FILLER_0_119_563 ();
 sg13g2_fill_2 FILLER_0_119_570 ();
 sg13g2_fill_1 FILLER_0_119_572 ();
 sg13g2_fill_2 FILLER_0_119_578 ();
 sg13g2_fill_1 FILLER_0_119_580 ();
 sg13g2_fill_2 FILLER_0_119_585 ();
 sg13g2_fill_2 FILLER_0_119_613 ();
 sg13g2_fill_2 FILLER_0_119_621 ();
 sg13g2_fill_8 FILLER_0_119_629 ();
 sg13g2_fill_4 FILLER_0_119_637 ();
 sg13g2_fill_2 FILLER_0_119_641 ();
 sg13g2_fill_1 FILLER_0_119_643 ();
 sg13g2_fill_2 FILLER_0_119_649 ();
 sg13g2_fill_4 FILLER_0_119_655 ();
 sg13g2_fill_1 FILLER_0_119_659 ();
 sg13g2_fill_4 FILLER_0_119_665 ();
 sg13g2_fill_1 FILLER_0_119_669 ();
 sg13g2_fill_2 FILLER_0_119_675 ();
 sg13g2_fill_4 FILLER_0_119_682 ();
 sg13g2_fill_1 FILLER_0_119_686 ();
 sg13g2_fill_2 FILLER_0_119_713 ();
 sg13g2_fill_8 FILLER_0_119_725 ();
 sg13g2_fill_4 FILLER_0_119_733 ();
 sg13g2_fill_2 FILLER_0_119_737 ();
 sg13g2_fill_1 FILLER_0_119_739 ();
 sg13g2_fill_4 FILLER_0_119_745 ();
 sg13g2_fill_1 FILLER_0_119_749 ();
 sg13g2_fill_4 FILLER_0_119_755 ();
 sg13g2_fill_2 FILLER_0_119_759 ();
 sg13g2_fill_2 FILLER_0_119_787 ();
 sg13g2_fill_8 FILLER_0_119_794 ();
 sg13g2_fill_8 FILLER_0_119_802 ();
 sg13g2_fill_4 FILLER_0_119_815 ();
 sg13g2_fill_2 FILLER_0_119_819 ();
 sg13g2_fill_2 FILLER_0_119_826 ();
 sg13g2_fill_2 FILLER_0_119_833 ();
 sg13g2_fill_4 FILLER_0_119_839 ();
 sg13g2_fill_1 FILLER_0_119_843 ();
 sg13g2_fill_8 FILLER_0_119_848 ();
 sg13g2_fill_8 FILLER_0_119_856 ();
 sg13g2_fill_2 FILLER_0_119_890 ();
 sg13g2_fill_8 FILLER_0_119_897 ();
 sg13g2_fill_8 FILLER_0_119_905 ();
 sg13g2_fill_8 FILLER_0_119_913 ();
 sg13g2_fill_4 FILLER_0_119_921 ();
 sg13g2_fill_2 FILLER_0_119_925 ();
 sg13g2_fill_8 FILLER_0_119_931 ();
 sg13g2_fill_2 FILLER_0_119_939 ();
 sg13g2_fill_1 FILLER_0_119_941 ();
 sg13g2_fill_2 FILLER_0_119_946 ();
 sg13g2_fill_1 FILLER_0_119_948 ();
 sg13g2_fill_2 FILLER_0_119_955 ();
 sg13g2_fill_2 FILLER_0_119_962 ();
 sg13g2_fill_2 FILLER_0_119_969 ();
 sg13g2_fill_8 FILLER_0_119_975 ();
 sg13g2_fill_8 FILLER_0_119_983 ();
 sg13g2_fill_4 FILLER_0_119_991 ();
 sg13g2_fill_2 FILLER_0_119_995 ();
 sg13g2_fill_1 FILLER_0_119_997 ();
 sg13g2_fill_8 FILLER_0_119_1003 ();
 sg13g2_fill_4 FILLER_0_119_1011 ();
 sg13g2_fill_2 FILLER_0_119_1020 ();
 sg13g2_fill_1 FILLER_0_119_1022 ();
 sg13g2_fill_4 FILLER_0_119_1028 ();
 sg13g2_fill_4 FILLER_0_119_1038 ();
 sg13g2_fill_4 FILLER_0_119_1046 ();
 sg13g2_fill_1 FILLER_0_119_1050 ();
 sg13g2_fill_2 FILLER_0_119_1057 ();
 sg13g2_fill_2 FILLER_0_119_1063 ();
 sg13g2_fill_1 FILLER_0_119_1065 ();
 sg13g2_fill_8 FILLER_0_119_1073 ();
 sg13g2_fill_8 FILLER_0_119_1081 ();
 sg13g2_fill_8 FILLER_0_119_1089 ();
 sg13g2_fill_8 FILLER_0_119_1097 ();
 sg13g2_fill_8 FILLER_0_119_1105 ();
 sg13g2_fill_8 FILLER_0_119_1113 ();
 sg13g2_fill_8 FILLER_0_119_1121 ();
 sg13g2_fill_8 FILLER_0_119_1129 ();
 sg13g2_fill_8 FILLER_0_119_1137 ();
 sg13g2_fill_8 FILLER_0_119_1145 ();
 sg13g2_fill_2 FILLER_0_119_1153 ();
 sg13g2_fill_8 FILLER_0_119_1159 ();
 sg13g2_fill_8 FILLER_0_119_1167 ();
 sg13g2_fill_8 FILLER_0_119_1175 ();
 sg13g2_fill_2 FILLER_0_119_1183 ();
 sg13g2_fill_8 FILLER_0_119_1189 ();
 sg13g2_fill_8 FILLER_0_119_1197 ();
 sg13g2_fill_4 FILLER_0_119_1205 ();
 sg13g2_fill_2 FILLER_0_119_1217 ();
 sg13g2_fill_1 FILLER_0_119_1219 ();
 sg13g2_fill_2 FILLER_0_119_1228 ();
 sg13g2_fill_1 FILLER_0_119_1230 ();
 sg13g2_fill_2 FILLER_0_119_1236 ();
 sg13g2_fill_1 FILLER_0_119_1238 ();
 sg13g2_fill_2 FILLER_0_119_1247 ();
 sg13g2_fill_1 FILLER_0_119_1249 ();
 sg13g2_fill_4 FILLER_0_119_1260 ();
 sg13g2_fill_2 FILLER_0_119_1264 ();
 sg13g2_fill_2 FILLER_0_119_1274 ();
 sg13g2_fill_2 FILLER_0_119_1280 ();
 sg13g2_fill_1 FILLER_0_119_1282 ();
 sg13g2_fill_4 FILLER_0_119_1286 ();
 sg13g2_fill_2 FILLER_0_119_1290 ();
 sg13g2_fill_1 FILLER_0_119_1296 ();
 sg13g2_fill_8 FILLER_0_120_0 ();
 sg13g2_fill_8 FILLER_0_120_8 ();
 sg13g2_fill_8 FILLER_0_120_16 ();
 sg13g2_fill_8 FILLER_0_120_24 ();
 sg13g2_fill_8 FILLER_0_120_32 ();
 sg13g2_fill_8 FILLER_0_120_40 ();
 sg13g2_fill_8 FILLER_0_120_48 ();
 sg13g2_fill_8 FILLER_0_120_56 ();
 sg13g2_fill_8 FILLER_0_120_64 ();
 sg13g2_fill_8 FILLER_0_120_72 ();
 sg13g2_fill_8 FILLER_0_120_80 ();
 sg13g2_fill_8 FILLER_0_120_88 ();
 sg13g2_fill_8 FILLER_0_120_96 ();
 sg13g2_fill_8 FILLER_0_120_104 ();
 sg13g2_fill_8 FILLER_0_120_112 ();
 sg13g2_fill_8 FILLER_0_120_120 ();
 sg13g2_fill_8 FILLER_0_120_128 ();
 sg13g2_fill_8 FILLER_0_120_136 ();
 sg13g2_fill_8 FILLER_0_120_144 ();
 sg13g2_fill_8 FILLER_0_120_152 ();
 sg13g2_fill_8 FILLER_0_120_160 ();
 sg13g2_fill_8 FILLER_0_120_168 ();
 sg13g2_fill_8 FILLER_0_120_176 ();
 sg13g2_fill_8 FILLER_0_120_184 ();
 sg13g2_fill_8 FILLER_0_120_192 ();
 sg13g2_fill_8 FILLER_0_120_200 ();
 sg13g2_fill_8 FILLER_0_120_208 ();
 sg13g2_fill_8 FILLER_0_120_216 ();
 sg13g2_fill_8 FILLER_0_120_224 ();
 sg13g2_fill_8 FILLER_0_120_232 ();
 sg13g2_fill_4 FILLER_0_120_261 ();
 sg13g2_fill_4 FILLER_0_120_270 ();
 sg13g2_fill_1 FILLER_0_120_274 ();
 sg13g2_fill_8 FILLER_0_120_279 ();
 sg13g2_fill_1 FILLER_0_120_287 ();
 sg13g2_fill_4 FILLER_0_120_298 ();
 sg13g2_fill_1 FILLER_0_120_302 ();
 sg13g2_fill_2 FILLER_0_120_308 ();
 sg13g2_fill_8 FILLER_0_120_315 ();
 sg13g2_fill_8 FILLER_0_120_323 ();
 sg13g2_fill_8 FILLER_0_120_331 ();
 sg13g2_fill_8 FILLER_0_120_339 ();
 sg13g2_fill_8 FILLER_0_120_347 ();
 sg13g2_fill_8 FILLER_0_120_355 ();
 sg13g2_fill_1 FILLER_0_120_363 ();
 sg13g2_fill_8 FILLER_0_120_368 ();
 sg13g2_fill_8 FILLER_0_120_376 ();
 sg13g2_fill_4 FILLER_0_120_384 ();
 sg13g2_fill_2 FILLER_0_120_392 ();
 sg13g2_fill_2 FILLER_0_120_399 ();
 sg13g2_fill_8 FILLER_0_120_411 ();
 sg13g2_fill_8 FILLER_0_120_419 ();
 sg13g2_fill_4 FILLER_0_120_427 ();
 sg13g2_fill_1 FILLER_0_120_431 ();
 sg13g2_fill_2 FILLER_0_120_438 ();
 sg13g2_fill_8 FILLER_0_120_445 ();
 sg13g2_fill_2 FILLER_0_120_453 ();
 sg13g2_fill_1 FILLER_0_120_455 ();
 sg13g2_fill_2 FILLER_0_120_461 ();
 sg13g2_fill_8 FILLER_0_120_467 ();
 sg13g2_fill_8 FILLER_0_120_475 ();
 sg13g2_fill_8 FILLER_0_120_483 ();
 sg13g2_fill_8 FILLER_0_120_491 ();
 sg13g2_fill_8 FILLER_0_120_499 ();
 sg13g2_fill_1 FILLER_0_120_507 ();
 sg13g2_fill_8 FILLER_0_120_534 ();
 sg13g2_fill_8 FILLER_0_120_546 ();
 sg13g2_fill_4 FILLER_0_120_554 ();
 sg13g2_fill_2 FILLER_0_120_558 ();
 sg13g2_fill_8 FILLER_0_120_565 ();
 sg13g2_fill_2 FILLER_0_120_573 ();
 sg13g2_fill_2 FILLER_0_120_601 ();
 sg13g2_fill_2 FILLER_0_120_608 ();
 sg13g2_fill_1 FILLER_0_120_610 ();
 sg13g2_fill_2 FILLER_0_120_616 ();
 sg13g2_fill_2 FILLER_0_120_624 ();
 sg13g2_fill_2 FILLER_0_120_635 ();
 sg13g2_fill_2 FILLER_0_120_641 ();
 sg13g2_fill_2 FILLER_0_120_648 ();
 sg13g2_fill_2 FILLER_0_120_676 ();
 sg13g2_fill_2 FILLER_0_120_682 ();
 sg13g2_fill_1 FILLER_0_120_684 ();
 sg13g2_fill_4 FILLER_0_120_690 ();
 sg13g2_fill_2 FILLER_0_120_694 ();
 sg13g2_fill_2 FILLER_0_120_700 ();
 sg13g2_fill_4 FILLER_0_120_710 ();
 sg13g2_fill_2 FILLER_0_120_714 ();
 sg13g2_fill_8 FILLER_0_120_721 ();
 sg13g2_fill_1 FILLER_0_120_729 ();
 sg13g2_fill_8 FILLER_0_120_735 ();
 sg13g2_fill_2 FILLER_0_120_743 ();
 sg13g2_fill_2 FILLER_0_120_750 ();
 sg13g2_fill_8 FILLER_0_120_756 ();
 sg13g2_fill_8 FILLER_0_120_764 ();
 sg13g2_fill_8 FILLER_0_120_772 ();
 sg13g2_fill_8 FILLER_0_120_780 ();
 sg13g2_fill_8 FILLER_0_120_788 ();
 sg13g2_fill_1 FILLER_0_120_796 ();
 sg13g2_fill_4 FILLER_0_120_807 ();
 sg13g2_fill_8 FILLER_0_120_816 ();
 sg13g2_fill_8 FILLER_0_120_824 ();
 sg13g2_fill_8 FILLER_0_120_832 ();
 sg13g2_fill_1 FILLER_0_120_840 ();
 sg13g2_fill_2 FILLER_0_120_845 ();
 sg13g2_fill_8 FILLER_0_120_857 ();
 sg13g2_fill_8 FILLER_0_120_865 ();
 sg13g2_fill_4 FILLER_0_120_873 ();
 sg13g2_fill_8 FILLER_0_120_883 ();
 sg13g2_fill_8 FILLER_0_120_891 ();
 sg13g2_fill_1 FILLER_0_120_899 ();
 sg13g2_fill_8 FILLER_0_120_926 ();
 sg13g2_fill_8 FILLER_0_120_934 ();
 sg13g2_fill_8 FILLER_0_120_942 ();
 sg13g2_fill_8 FILLER_0_120_950 ();
 sg13g2_fill_4 FILLER_0_120_958 ();
 sg13g2_fill_2 FILLER_0_120_962 ();
 sg13g2_fill_8 FILLER_0_120_967 ();
 sg13g2_fill_8 FILLER_0_120_975 ();
 sg13g2_fill_4 FILLER_0_120_983 ();
 sg13g2_fill_2 FILLER_0_120_987 ();
 sg13g2_fill_1 FILLER_0_120_989 ();
 sg13g2_fill_8 FILLER_0_120_996 ();
 sg13g2_fill_8 FILLER_0_120_1004 ();
 sg13g2_fill_8 FILLER_0_120_1012 ();
 sg13g2_fill_4 FILLER_0_120_1020 ();
 sg13g2_fill_2 FILLER_0_120_1024 ();
 sg13g2_fill_8 FILLER_0_120_1031 ();
 sg13g2_fill_1 FILLER_0_120_1039 ();
 sg13g2_fill_2 FILLER_0_120_1046 ();
 sg13g2_fill_1 FILLER_0_120_1048 ();
 sg13g2_fill_2 FILLER_0_120_1053 ();
 sg13g2_fill_2 FILLER_0_120_1060 ();
 sg13g2_fill_4 FILLER_0_120_1066 ();
 sg13g2_fill_8 FILLER_0_120_1075 ();
 sg13g2_fill_4 FILLER_0_120_1083 ();
 sg13g2_fill_8 FILLER_0_120_1092 ();
 sg13g2_fill_2 FILLER_0_120_1100 ();
 sg13g2_fill_2 FILLER_0_120_1107 ();
 sg13g2_fill_4 FILLER_0_120_1114 ();
 sg13g2_fill_2 FILLER_0_120_1118 ();
 sg13g2_fill_1 FILLER_0_120_1120 ();
 sg13g2_fill_8 FILLER_0_120_1131 ();
 sg13g2_fill_8 FILLER_0_120_1139 ();
 sg13g2_fill_8 FILLER_0_120_1147 ();
 sg13g2_fill_8 FILLER_0_120_1155 ();
 sg13g2_fill_8 FILLER_0_120_1163 ();
 sg13g2_fill_8 FILLER_0_120_1171 ();
 sg13g2_fill_8 FILLER_0_120_1179 ();
 sg13g2_fill_8 FILLER_0_120_1187 ();
 sg13g2_fill_8 FILLER_0_120_1195 ();
 sg13g2_fill_8 FILLER_0_120_1203 ();
 sg13g2_fill_8 FILLER_0_120_1211 ();
 sg13g2_fill_4 FILLER_0_120_1219 ();
 sg13g2_fill_2 FILLER_0_120_1228 ();
 sg13g2_fill_2 FILLER_0_120_1235 ();
 sg13g2_fill_1 FILLER_0_120_1237 ();
 sg13g2_fill_2 FILLER_0_120_1246 ();
 sg13g2_fill_1 FILLER_0_120_1248 ();
 sg13g2_fill_2 FILLER_0_120_1259 ();
 sg13g2_fill_4 FILLER_0_120_1267 ();
 sg13g2_fill_1 FILLER_0_120_1271 ();
 sg13g2_fill_2 FILLER_0_120_1277 ();
 sg13g2_fill_2 FILLER_0_120_1283 ();
 sg13g2_fill_1 FILLER_0_120_1285 ();
 sg13g2_fill_4 FILLER_0_120_1290 ();
 sg13g2_fill_2 FILLER_0_120_1294 ();
 sg13g2_fill_1 FILLER_0_120_1296 ();
 sg13g2_fill_8 FILLER_0_121_0 ();
 sg13g2_fill_8 FILLER_0_121_8 ();
 sg13g2_fill_8 FILLER_0_121_16 ();
 sg13g2_fill_8 FILLER_0_121_24 ();
 sg13g2_fill_8 FILLER_0_121_32 ();
 sg13g2_fill_8 FILLER_0_121_40 ();
 sg13g2_fill_8 FILLER_0_121_48 ();
 sg13g2_fill_8 FILLER_0_121_56 ();
 sg13g2_fill_8 FILLER_0_121_64 ();
 sg13g2_fill_8 FILLER_0_121_72 ();
 sg13g2_fill_8 FILLER_0_121_80 ();
 sg13g2_fill_8 FILLER_0_121_88 ();
 sg13g2_fill_8 FILLER_0_121_96 ();
 sg13g2_fill_8 FILLER_0_121_104 ();
 sg13g2_fill_8 FILLER_0_121_112 ();
 sg13g2_fill_8 FILLER_0_121_120 ();
 sg13g2_fill_8 FILLER_0_121_128 ();
 sg13g2_fill_8 FILLER_0_121_136 ();
 sg13g2_fill_8 FILLER_0_121_144 ();
 sg13g2_fill_8 FILLER_0_121_152 ();
 sg13g2_fill_8 FILLER_0_121_160 ();
 sg13g2_fill_8 FILLER_0_121_168 ();
 sg13g2_fill_8 FILLER_0_121_176 ();
 sg13g2_fill_8 FILLER_0_121_184 ();
 sg13g2_fill_8 FILLER_0_121_192 ();
 sg13g2_fill_8 FILLER_0_121_200 ();
 sg13g2_fill_4 FILLER_0_121_208 ();
 sg13g2_fill_2 FILLER_0_121_212 ();
 sg13g2_fill_1 FILLER_0_121_214 ();
 sg13g2_fill_2 FILLER_0_121_241 ();
 sg13g2_fill_2 FILLER_0_121_269 ();
 sg13g2_fill_4 FILLER_0_121_276 ();
 sg13g2_fill_2 FILLER_0_121_280 ();
 sg13g2_fill_4 FILLER_0_121_287 ();
 sg13g2_fill_4 FILLER_0_121_295 ();
 sg13g2_fill_2 FILLER_0_121_299 ();
 sg13g2_fill_1 FILLER_0_121_301 ();
 sg13g2_fill_8 FILLER_0_121_328 ();
 sg13g2_fill_1 FILLER_0_121_336 ();
 sg13g2_fill_2 FILLER_0_121_363 ();
 sg13g2_fill_4 FILLER_0_121_370 ();
 sg13g2_fill_8 FILLER_0_121_378 ();
 sg13g2_fill_8 FILLER_0_121_386 ();
 sg13g2_fill_8 FILLER_0_121_394 ();
 sg13g2_fill_4 FILLER_0_121_402 ();
 sg13g2_fill_2 FILLER_0_121_406 ();
 sg13g2_fill_1 FILLER_0_121_408 ();
 sg13g2_fill_2 FILLER_0_121_413 ();
 sg13g2_fill_2 FILLER_0_121_420 ();
 sg13g2_fill_2 FILLER_0_121_429 ();
 sg13g2_fill_8 FILLER_0_121_436 ();
 sg13g2_fill_8 FILLER_0_121_444 ();
 sg13g2_fill_1 FILLER_0_121_452 ();
 sg13g2_fill_4 FILLER_0_121_479 ();
 sg13g2_fill_4 FILLER_0_121_504 ();
 sg13g2_fill_2 FILLER_0_121_513 ();
 sg13g2_fill_2 FILLER_0_121_541 ();
 sg13g2_fill_2 FILLER_0_121_553 ();
 sg13g2_fill_8 FILLER_0_121_560 ();
 sg13g2_fill_8 FILLER_0_121_568 ();
 sg13g2_fill_8 FILLER_0_121_576 ();
 sg13g2_fill_8 FILLER_0_121_584 ();
 sg13g2_fill_8 FILLER_0_121_592 ();
 sg13g2_fill_2 FILLER_0_121_610 ();
 sg13g2_fill_1 FILLER_0_121_612 ();
 sg13g2_fill_8 FILLER_0_121_617 ();
 sg13g2_fill_2 FILLER_0_121_625 ();
 sg13g2_fill_2 FILLER_0_121_632 ();
 sg13g2_fill_2 FILLER_0_121_639 ();
 sg13g2_fill_4 FILLER_0_121_646 ();
 sg13g2_fill_4 FILLER_0_121_655 ();
 sg13g2_fill_8 FILLER_0_121_663 ();
 sg13g2_fill_8 FILLER_0_121_671 ();
 sg13g2_fill_8 FILLER_0_121_679 ();
 sg13g2_fill_8 FILLER_0_121_687 ();
 sg13g2_fill_8 FILLER_0_121_695 ();
 sg13g2_fill_8 FILLER_0_121_703 ();
 sg13g2_fill_4 FILLER_0_121_711 ();
 sg13g2_fill_1 FILLER_0_121_715 ();
 sg13g2_fill_8 FILLER_0_121_742 ();
 sg13g2_fill_8 FILLER_0_121_750 ();
 sg13g2_fill_8 FILLER_0_121_758 ();
 sg13g2_fill_8 FILLER_0_121_766 ();
 sg13g2_fill_8 FILLER_0_121_774 ();
 sg13g2_fill_4 FILLER_0_121_782 ();
 sg13g2_fill_1 FILLER_0_121_786 ();
 sg13g2_fill_8 FILLER_0_121_813 ();
 sg13g2_fill_4 FILLER_0_121_821 ();
 sg13g2_fill_2 FILLER_0_121_825 ();
 sg13g2_fill_1 FILLER_0_121_827 ();
 sg13g2_fill_2 FILLER_0_121_833 ();
 sg13g2_fill_1 FILLER_0_121_835 ();
 sg13g2_fill_2 FILLER_0_121_862 ();
 sg13g2_fill_8 FILLER_0_121_869 ();
 sg13g2_fill_8 FILLER_0_121_877 ();
 sg13g2_fill_8 FILLER_0_121_885 ();
 sg13g2_fill_4 FILLER_0_121_893 ();
 sg13g2_fill_2 FILLER_0_121_897 ();
 sg13g2_fill_2 FILLER_0_121_904 ();
 sg13g2_fill_1 FILLER_0_121_906 ();
 sg13g2_fill_4 FILLER_0_121_911 ();
 sg13g2_fill_2 FILLER_0_121_915 ();
 sg13g2_fill_2 FILLER_0_121_921 ();
 sg13g2_fill_8 FILLER_0_121_928 ();
 sg13g2_fill_8 FILLER_0_121_936 ();
 sg13g2_fill_8 FILLER_0_121_944 ();
 sg13g2_fill_8 FILLER_0_121_952 ();
 sg13g2_fill_4 FILLER_0_121_960 ();
 sg13g2_fill_1 FILLER_0_121_964 ();
 sg13g2_fill_2 FILLER_0_121_972 ();
 sg13g2_fill_8 FILLER_0_121_980 ();
 sg13g2_fill_8 FILLER_0_121_988 ();
 sg13g2_fill_4 FILLER_0_121_996 ();
 sg13g2_fill_2 FILLER_0_121_1005 ();
 sg13g2_fill_8 FILLER_0_121_1011 ();
 sg13g2_fill_8 FILLER_0_121_1019 ();
 sg13g2_fill_8 FILLER_0_121_1027 ();
 sg13g2_fill_8 FILLER_0_121_1035 ();
 sg13g2_fill_4 FILLER_0_121_1043 ();
 sg13g2_fill_2 FILLER_0_121_1047 ();
 sg13g2_fill_1 FILLER_0_121_1049 ();
 sg13g2_fill_8 FILLER_0_121_1056 ();
 sg13g2_fill_2 FILLER_0_121_1064 ();
 sg13g2_fill_1 FILLER_0_121_1066 ();
 sg13g2_fill_8 FILLER_0_121_1075 ();
 sg13g2_fill_8 FILLER_0_121_1083 ();
 sg13g2_fill_8 FILLER_0_121_1091 ();
 sg13g2_fill_8 FILLER_0_121_1099 ();
 sg13g2_fill_8 FILLER_0_121_1107 ();
 sg13g2_fill_8 FILLER_0_121_1115 ();
 sg13g2_fill_8 FILLER_0_121_1127 ();
 sg13g2_fill_8 FILLER_0_121_1135 ();
 sg13g2_fill_8 FILLER_0_121_1143 ();
 sg13g2_fill_8 FILLER_0_121_1151 ();
 sg13g2_fill_8 FILLER_0_121_1159 ();
 sg13g2_fill_8 FILLER_0_121_1167 ();
 sg13g2_fill_8 FILLER_0_121_1175 ();
 sg13g2_fill_8 FILLER_0_121_1183 ();
 sg13g2_fill_1 FILLER_0_121_1191 ();
 sg13g2_fill_8 FILLER_0_121_1197 ();
 sg13g2_fill_8 FILLER_0_121_1205 ();
 sg13g2_fill_8 FILLER_0_121_1213 ();
 sg13g2_fill_2 FILLER_0_121_1221 ();
 sg13g2_fill_1 FILLER_0_121_1223 ();
 sg13g2_fill_2 FILLER_0_121_1227 ();
 sg13g2_fill_8 FILLER_0_121_1234 ();
 sg13g2_fill_8 FILLER_0_121_1242 ();
 sg13g2_fill_2 FILLER_0_121_1276 ();
 sg13g2_fill_2 FILLER_0_121_1282 ();
 sg13g2_fill_1 FILLER_0_121_1284 ();
 sg13g2_fill_8 FILLER_0_121_1289 ();
 sg13g2_fill_8 FILLER_0_122_0 ();
 sg13g2_fill_8 FILLER_0_122_8 ();
 sg13g2_fill_8 FILLER_0_122_16 ();
 sg13g2_fill_8 FILLER_0_122_24 ();
 sg13g2_fill_8 FILLER_0_122_32 ();
 sg13g2_fill_8 FILLER_0_122_40 ();
 sg13g2_fill_8 FILLER_0_122_48 ();
 sg13g2_fill_8 FILLER_0_122_56 ();
 sg13g2_fill_8 FILLER_0_122_64 ();
 sg13g2_fill_8 FILLER_0_122_72 ();
 sg13g2_fill_8 FILLER_0_122_80 ();
 sg13g2_fill_8 FILLER_0_122_88 ();
 sg13g2_fill_8 FILLER_0_122_96 ();
 sg13g2_fill_8 FILLER_0_122_104 ();
 sg13g2_fill_8 FILLER_0_122_112 ();
 sg13g2_fill_8 FILLER_0_122_120 ();
 sg13g2_fill_8 FILLER_0_122_128 ();
 sg13g2_fill_8 FILLER_0_122_136 ();
 sg13g2_fill_8 FILLER_0_122_144 ();
 sg13g2_fill_8 FILLER_0_122_152 ();
 sg13g2_fill_8 FILLER_0_122_160 ();
 sg13g2_fill_8 FILLER_0_122_168 ();
 sg13g2_fill_8 FILLER_0_122_176 ();
 sg13g2_fill_8 FILLER_0_122_184 ();
 sg13g2_fill_8 FILLER_0_122_192 ();
 sg13g2_fill_8 FILLER_0_122_200 ();
 sg13g2_fill_8 FILLER_0_122_208 ();
 sg13g2_fill_4 FILLER_0_122_216 ();
 sg13g2_fill_2 FILLER_0_122_220 ();
 sg13g2_fill_2 FILLER_0_122_227 ();
 sg13g2_fill_4 FILLER_0_122_233 ();
 sg13g2_fill_8 FILLER_0_122_242 ();
 sg13g2_fill_4 FILLER_0_122_250 ();
 sg13g2_fill_2 FILLER_0_122_254 ();
 sg13g2_fill_1 FILLER_0_122_256 ();
 sg13g2_fill_4 FILLER_0_122_263 ();
 sg13g2_fill_4 FILLER_0_122_293 ();
 sg13g2_fill_2 FILLER_0_122_297 ();
 sg13g2_fill_1 FILLER_0_122_299 ();
 sg13g2_fill_8 FILLER_0_122_305 ();
 sg13g2_fill_8 FILLER_0_122_313 ();
 sg13g2_fill_8 FILLER_0_122_321 ();
 sg13g2_fill_8 FILLER_0_122_329 ();
 sg13g2_fill_8 FILLER_0_122_337 ();
 sg13g2_fill_4 FILLER_0_122_345 ();
 sg13g2_fill_2 FILLER_0_122_349 ();
 sg13g2_fill_4 FILLER_0_122_356 ();
 sg13g2_fill_2 FILLER_0_122_360 ();
 sg13g2_fill_2 FILLER_0_122_383 ();
 sg13g2_fill_2 FILLER_0_122_406 ();
 sg13g2_fill_1 FILLER_0_122_408 ();
 sg13g2_fill_2 FILLER_0_122_414 ();
 sg13g2_fill_8 FILLER_0_122_442 ();
 sg13g2_fill_8 FILLER_0_122_450 ();
 sg13g2_fill_4 FILLER_0_122_458 ();
 sg13g2_fill_2 FILLER_0_122_467 ();
 sg13g2_fill_4 FILLER_0_122_495 ();
 sg13g2_fill_4 FILLER_0_122_508 ();
 sg13g2_fill_2 FILLER_0_122_512 ();
 sg13g2_fill_4 FILLER_0_122_519 ();
 sg13g2_fill_8 FILLER_0_122_527 ();
 sg13g2_fill_8 FILLER_0_122_535 ();
 sg13g2_fill_2 FILLER_0_122_543 ();
 sg13g2_fill_2 FILLER_0_122_550 ();
 sg13g2_fill_2 FILLER_0_122_557 ();
 sg13g2_fill_4 FILLER_0_122_565 ();
 sg13g2_fill_8 FILLER_0_122_574 ();
 sg13g2_fill_8 FILLER_0_122_582 ();
 sg13g2_fill_8 FILLER_0_122_590 ();
 sg13g2_fill_8 FILLER_0_122_598 ();
 sg13g2_fill_2 FILLER_0_122_606 ();
 sg13g2_fill_1 FILLER_0_122_608 ();
 sg13g2_fill_2 FILLER_0_122_614 ();
 sg13g2_fill_8 FILLER_0_122_628 ();
 sg13g2_fill_8 FILLER_0_122_636 ();
 sg13g2_fill_8 FILLER_0_122_644 ();
 sg13g2_fill_8 FILLER_0_122_652 ();
 sg13g2_fill_8 FILLER_0_122_660 ();
 sg13g2_fill_8 FILLER_0_122_668 ();
 sg13g2_fill_8 FILLER_0_122_676 ();
 sg13g2_fill_8 FILLER_0_122_684 ();
 sg13g2_fill_8 FILLER_0_122_692 ();
 sg13g2_fill_1 FILLER_0_122_700 ();
 sg13g2_fill_4 FILLER_0_122_706 ();
 sg13g2_fill_2 FILLER_0_122_714 ();
 sg13g2_fill_1 FILLER_0_122_716 ();
 sg13g2_fill_8 FILLER_0_122_722 ();
 sg13g2_fill_8 FILLER_0_122_730 ();
 sg13g2_fill_8 FILLER_0_122_738 ();
 sg13g2_fill_8 FILLER_0_122_746 ();
 sg13g2_fill_8 FILLER_0_122_754 ();
 sg13g2_fill_8 FILLER_0_122_762 ();
 sg13g2_fill_8 FILLER_0_122_770 ();
 sg13g2_fill_8 FILLER_0_122_778 ();
 sg13g2_fill_2 FILLER_0_122_790 ();
 sg13g2_fill_2 FILLER_0_122_797 ();
 sg13g2_fill_2 FILLER_0_122_803 ();
 sg13g2_fill_1 FILLER_0_122_805 ();
 sg13g2_fill_8 FILLER_0_122_810 ();
 sg13g2_fill_8 FILLER_0_122_818 ();
 sg13g2_fill_8 FILLER_0_122_826 ();
 sg13g2_fill_4 FILLER_0_122_834 ();
 sg13g2_fill_1 FILLER_0_122_838 ();
 sg13g2_fill_2 FILLER_0_122_844 ();
 sg13g2_fill_8 FILLER_0_122_850 ();
 sg13g2_fill_8 FILLER_0_122_858 ();
 sg13g2_fill_2 FILLER_0_122_866 ();
 sg13g2_fill_1 FILLER_0_122_868 ();
 sg13g2_fill_2 FILLER_0_122_895 ();
 sg13g2_fill_8 FILLER_0_122_902 ();
 sg13g2_fill_8 FILLER_0_122_910 ();
 sg13g2_fill_4 FILLER_0_122_926 ();
 sg13g2_fill_1 FILLER_0_122_930 ();
 sg13g2_fill_8 FILLER_0_122_936 ();
 sg13g2_fill_8 FILLER_0_122_944 ();
 sg13g2_fill_8 FILLER_0_122_952 ();
 sg13g2_fill_8 FILLER_0_122_960 ();
 sg13g2_fill_4 FILLER_0_122_968 ();
 sg13g2_fill_2 FILLER_0_122_977 ();
 sg13g2_fill_2 FILLER_0_122_987 ();
 sg13g2_fill_1 FILLER_0_122_989 ();
 sg13g2_fill_2 FILLER_0_122_995 ();
 sg13g2_fill_2 FILLER_0_122_1003 ();
 sg13g2_fill_8 FILLER_0_122_1010 ();
 sg13g2_fill_8 FILLER_0_122_1018 ();
 sg13g2_fill_8 FILLER_0_122_1026 ();
 sg13g2_fill_4 FILLER_0_122_1034 ();
 sg13g2_fill_2 FILLER_0_122_1038 ();
 sg13g2_fill_8 FILLER_0_122_1045 ();
 sg13g2_fill_2 FILLER_0_122_1061 ();
 sg13g2_fill_8 FILLER_0_122_1068 ();
 sg13g2_fill_2 FILLER_0_122_1076 ();
 sg13g2_fill_8 FILLER_0_122_1081 ();
 sg13g2_fill_4 FILLER_0_122_1089 ();
 sg13g2_fill_2 FILLER_0_122_1093 ();
 sg13g2_fill_1 FILLER_0_122_1095 ();
 sg13g2_fill_2 FILLER_0_122_1101 ();
 sg13g2_fill_2 FILLER_0_122_1109 ();
 sg13g2_fill_4 FILLER_0_122_1118 ();
 sg13g2_fill_2 FILLER_0_122_1127 ();
 sg13g2_fill_4 FILLER_0_122_1136 ();
 sg13g2_fill_8 FILLER_0_122_1145 ();
 sg13g2_fill_8 FILLER_0_122_1153 ();
 sg13g2_fill_4 FILLER_0_122_1161 ();
 sg13g2_fill_2 FILLER_0_122_1165 ();
 sg13g2_fill_4 FILLER_0_122_1171 ();
 sg13g2_fill_2 FILLER_0_122_1175 ();
 sg13g2_fill_1 FILLER_0_122_1177 ();
 sg13g2_fill_4 FILLER_0_122_1186 ();
 sg13g2_fill_1 FILLER_0_122_1190 ();
 sg13g2_fill_4 FILLER_0_122_1199 ();
 sg13g2_fill_1 FILLER_0_122_1203 ();
 sg13g2_fill_2 FILLER_0_122_1212 ();
 sg13g2_fill_8 FILLER_0_122_1218 ();
 sg13g2_fill_8 FILLER_0_122_1231 ();
 sg13g2_fill_8 FILLER_0_122_1239 ();
 sg13g2_fill_8 FILLER_0_122_1247 ();
 sg13g2_fill_8 FILLER_0_122_1255 ();
 sg13g2_fill_2 FILLER_0_122_1263 ();
 sg13g2_fill_8 FILLER_0_122_1269 ();
 sg13g2_fill_4 FILLER_0_122_1277 ();
 sg13g2_fill_2 FILLER_0_122_1281 ();
 sg13g2_fill_8 FILLER_0_122_1287 ();
 sg13g2_fill_2 FILLER_0_122_1295 ();
 sg13g2_fill_8 FILLER_0_123_0 ();
 sg13g2_fill_8 FILLER_0_123_8 ();
 sg13g2_fill_8 FILLER_0_123_16 ();
 sg13g2_fill_8 FILLER_0_123_24 ();
 sg13g2_fill_8 FILLER_0_123_32 ();
 sg13g2_fill_8 FILLER_0_123_40 ();
 sg13g2_fill_8 FILLER_0_123_48 ();
 sg13g2_fill_8 FILLER_0_123_56 ();
 sg13g2_fill_8 FILLER_0_123_64 ();
 sg13g2_fill_8 FILLER_0_123_72 ();
 sg13g2_fill_8 FILLER_0_123_80 ();
 sg13g2_fill_8 FILLER_0_123_88 ();
 sg13g2_fill_8 FILLER_0_123_96 ();
 sg13g2_fill_8 FILLER_0_123_104 ();
 sg13g2_fill_8 FILLER_0_123_112 ();
 sg13g2_fill_8 FILLER_0_123_120 ();
 sg13g2_fill_8 FILLER_0_123_128 ();
 sg13g2_fill_8 FILLER_0_123_136 ();
 sg13g2_fill_8 FILLER_0_123_144 ();
 sg13g2_fill_8 FILLER_0_123_152 ();
 sg13g2_fill_8 FILLER_0_123_160 ();
 sg13g2_fill_8 FILLER_0_123_168 ();
 sg13g2_fill_8 FILLER_0_123_176 ();
 sg13g2_fill_8 FILLER_0_123_184 ();
 sg13g2_fill_8 FILLER_0_123_192 ();
 sg13g2_fill_8 FILLER_0_123_200 ();
 sg13g2_fill_8 FILLER_0_123_208 ();
 sg13g2_fill_8 FILLER_0_123_216 ();
 sg13g2_fill_8 FILLER_0_123_224 ();
 sg13g2_fill_8 FILLER_0_123_232 ();
 sg13g2_fill_4 FILLER_0_123_240 ();
 sg13g2_fill_1 FILLER_0_123_244 ();
 sg13g2_fill_2 FILLER_0_123_250 ();
 sg13g2_fill_8 FILLER_0_123_256 ();
 sg13g2_fill_8 FILLER_0_123_264 ();
 sg13g2_fill_4 FILLER_0_123_272 ();
 sg13g2_fill_2 FILLER_0_123_276 ();
 sg13g2_fill_1 FILLER_0_123_278 ();
 sg13g2_fill_4 FILLER_0_123_284 ();
 sg13g2_fill_8 FILLER_0_123_292 ();
 sg13g2_fill_8 FILLER_0_123_300 ();
 sg13g2_fill_8 FILLER_0_123_308 ();
 sg13g2_fill_8 FILLER_0_123_316 ();
 sg13g2_fill_8 FILLER_0_123_324 ();
 sg13g2_fill_8 FILLER_0_123_332 ();
 sg13g2_fill_4 FILLER_0_123_340 ();
 sg13g2_fill_2 FILLER_0_123_344 ();
 sg13g2_fill_2 FILLER_0_123_372 ();
 sg13g2_fill_2 FILLER_0_123_378 ();
 sg13g2_fill_2 FILLER_0_123_390 ();
 sg13g2_fill_2 FILLER_0_123_397 ();
 sg13g2_fill_8 FILLER_0_123_425 ();
 sg13g2_fill_8 FILLER_0_123_433 ();
 sg13g2_fill_8 FILLER_0_123_467 ();
 sg13g2_fill_4 FILLER_0_123_475 ();
 sg13g2_fill_8 FILLER_0_123_483 ();
 sg13g2_fill_2 FILLER_0_123_491 ();
 sg13g2_fill_8 FILLER_0_123_498 ();
 sg13g2_fill_8 FILLER_0_123_506 ();
 sg13g2_fill_8 FILLER_0_123_514 ();
 sg13g2_fill_8 FILLER_0_123_522 ();
 sg13g2_fill_8 FILLER_0_123_530 ();
 sg13g2_fill_8 FILLER_0_123_538 ();
 sg13g2_fill_2 FILLER_0_123_546 ();
 sg13g2_fill_4 FILLER_0_123_552 ();
 sg13g2_fill_1 FILLER_0_123_556 ();
 sg13g2_fill_2 FILLER_0_123_561 ();
 sg13g2_fill_4 FILLER_0_123_589 ();
 sg13g2_fill_2 FILLER_0_123_593 ();
 sg13g2_fill_4 FILLER_0_123_616 ();
 sg13g2_fill_2 FILLER_0_123_620 ();
 sg13g2_fill_1 FILLER_0_123_622 ();
 sg13g2_fill_2 FILLER_0_123_631 ();
 sg13g2_fill_8 FILLER_0_123_637 ();
 sg13g2_fill_2 FILLER_0_123_645 ();
 sg13g2_fill_2 FILLER_0_123_652 ();
 sg13g2_fill_2 FILLER_0_123_658 ();
 sg13g2_fill_8 FILLER_0_123_681 ();
 sg13g2_fill_4 FILLER_0_123_689 ();
 sg13g2_fill_2 FILLER_0_123_719 ();
 sg13g2_fill_4 FILLER_0_123_725 ();
 sg13g2_fill_2 FILLER_0_123_729 ();
 sg13g2_fill_2 FILLER_0_123_736 ();
 sg13g2_fill_1 FILLER_0_123_738 ();
 sg13g2_fill_2 FILLER_0_123_765 ();
 sg13g2_fill_8 FILLER_0_123_772 ();
 sg13g2_fill_8 FILLER_0_123_786 ();
 sg13g2_fill_8 FILLER_0_123_794 ();
 sg13g2_fill_2 FILLER_0_123_802 ();
 sg13g2_fill_1 FILLER_0_123_804 ();
 sg13g2_fill_2 FILLER_0_123_810 ();
 sg13g2_fill_4 FILLER_0_123_818 ();
 sg13g2_fill_2 FILLER_0_123_822 ();
 sg13g2_fill_1 FILLER_0_123_824 ();
 sg13g2_fill_4 FILLER_0_123_830 ();
 sg13g2_fill_8 FILLER_0_123_838 ();
 sg13g2_fill_4 FILLER_0_123_846 ();
 sg13g2_fill_2 FILLER_0_123_850 ();
 sg13g2_fill_2 FILLER_0_123_856 ();
 sg13g2_fill_1 FILLER_0_123_858 ();
 sg13g2_fill_2 FILLER_0_123_885 ();
 sg13g2_fill_2 FILLER_0_123_897 ();
 sg13g2_fill_2 FILLER_0_123_904 ();
 sg13g2_fill_2 FILLER_0_123_932 ();
 sg13g2_fill_8 FILLER_0_123_939 ();
 sg13g2_fill_8 FILLER_0_123_947 ();
 sg13g2_fill_8 FILLER_0_123_955 ();
 sg13g2_fill_8 FILLER_0_123_963 ();
 sg13g2_fill_8 FILLER_0_123_971 ();
 sg13g2_fill_8 FILLER_0_123_979 ();
 sg13g2_fill_8 FILLER_0_123_987 ();
 sg13g2_fill_2 FILLER_0_123_999 ();
 sg13g2_fill_2 FILLER_0_123_1006 ();
 sg13g2_fill_2 FILLER_0_123_1014 ();
 sg13g2_fill_8 FILLER_0_123_1021 ();
 sg13g2_fill_2 FILLER_0_123_1029 ();
 sg13g2_fill_1 FILLER_0_123_1031 ();
 sg13g2_fill_2 FILLER_0_123_1053 ();
 sg13g2_fill_2 FILLER_0_123_1060 ();
 sg13g2_fill_1 FILLER_0_123_1062 ();
 sg13g2_fill_2 FILLER_0_123_1069 ();
 sg13g2_fill_2 FILLER_0_123_1076 ();
 sg13g2_fill_1 FILLER_0_123_1078 ();
 sg13g2_fill_2 FILLER_0_123_1083 ();
 sg13g2_fill_8 FILLER_0_123_1090 ();
 sg13g2_fill_4 FILLER_0_123_1098 ();
 sg13g2_fill_1 FILLER_0_123_1102 ();
 sg13g2_fill_2 FILLER_0_123_1108 ();
 sg13g2_fill_1 FILLER_0_123_1110 ();
 sg13g2_fill_2 FILLER_0_123_1121 ();
 sg13g2_fill_4 FILLER_0_123_1131 ();
 sg13g2_fill_4 FILLER_0_123_1139 ();
 sg13g2_fill_2 FILLER_0_123_1143 ();
 sg13g2_fill_1 FILLER_0_123_1145 ();
 sg13g2_fill_4 FILLER_0_123_1152 ();
 sg13g2_fill_1 FILLER_0_123_1156 ();
 sg13g2_fill_2 FILLER_0_123_1167 ();
 sg13g2_fill_8 FILLER_0_123_1179 ();
 sg13g2_fill_2 FILLER_0_123_1187 ();
 sg13g2_fill_2 FILLER_0_123_1193 ();
 sg13g2_fill_1 FILLER_0_123_1195 ();
 sg13g2_fill_2 FILLER_0_123_1201 ();
 sg13g2_fill_2 FILLER_0_123_1210 ();
 sg13g2_fill_1 FILLER_0_123_1212 ();
 sg13g2_fill_2 FILLER_0_123_1218 ();
 sg13g2_fill_1 FILLER_0_123_1220 ();
 sg13g2_fill_8 FILLER_0_123_1226 ();
 sg13g2_fill_8 FILLER_0_123_1234 ();
 sg13g2_fill_4 FILLER_0_123_1242 ();
 sg13g2_fill_2 FILLER_0_123_1251 ();
 sg13g2_fill_8 FILLER_0_123_1257 ();
 sg13g2_fill_8 FILLER_0_123_1265 ();
 sg13g2_fill_2 FILLER_0_123_1273 ();
 sg13g2_fill_1 FILLER_0_123_1275 ();
 sg13g2_fill_8 FILLER_0_123_1284 ();
 sg13g2_fill_1 FILLER_0_123_1296 ();
 sg13g2_fill_8 FILLER_0_124_0 ();
 sg13g2_fill_8 FILLER_0_124_8 ();
 sg13g2_fill_8 FILLER_0_124_16 ();
 sg13g2_fill_8 FILLER_0_124_24 ();
 sg13g2_fill_8 FILLER_0_124_32 ();
 sg13g2_fill_8 FILLER_0_124_40 ();
 sg13g2_fill_8 FILLER_0_124_48 ();
 sg13g2_fill_8 FILLER_0_124_56 ();
 sg13g2_fill_8 FILLER_0_124_64 ();
 sg13g2_fill_8 FILLER_0_124_72 ();
 sg13g2_fill_8 FILLER_0_124_80 ();
 sg13g2_fill_8 FILLER_0_124_88 ();
 sg13g2_fill_8 FILLER_0_124_96 ();
 sg13g2_fill_8 FILLER_0_124_104 ();
 sg13g2_fill_8 FILLER_0_124_112 ();
 sg13g2_fill_8 FILLER_0_124_120 ();
 sg13g2_fill_8 FILLER_0_124_128 ();
 sg13g2_fill_8 FILLER_0_124_136 ();
 sg13g2_fill_8 FILLER_0_124_144 ();
 sg13g2_fill_8 FILLER_0_124_152 ();
 sg13g2_fill_8 FILLER_0_124_160 ();
 sg13g2_fill_8 FILLER_0_124_168 ();
 sg13g2_fill_8 FILLER_0_124_176 ();
 sg13g2_fill_8 FILLER_0_124_184 ();
 sg13g2_fill_8 FILLER_0_124_192 ();
 sg13g2_fill_8 FILLER_0_124_200 ();
 sg13g2_fill_8 FILLER_0_124_208 ();
 sg13g2_fill_8 FILLER_0_124_216 ();
 sg13g2_fill_8 FILLER_0_124_224 ();
 sg13g2_fill_8 FILLER_0_124_232 ();
 sg13g2_fill_8 FILLER_0_124_240 ();
 sg13g2_fill_8 FILLER_0_124_248 ();
 sg13g2_fill_8 FILLER_0_124_256 ();
 sg13g2_fill_8 FILLER_0_124_264 ();
 sg13g2_fill_2 FILLER_0_124_272 ();
 sg13g2_fill_8 FILLER_0_124_300 ();
 sg13g2_fill_8 FILLER_0_124_308 ();
 sg13g2_fill_8 FILLER_0_124_316 ();
 sg13g2_fill_8 FILLER_0_124_324 ();
 sg13g2_fill_4 FILLER_0_124_332 ();
 sg13g2_fill_8 FILLER_0_124_341 ();
 sg13g2_fill_8 FILLER_0_124_349 ();
 sg13g2_fill_8 FILLER_0_124_357 ();
 sg13g2_fill_1 FILLER_0_124_365 ();
 sg13g2_fill_8 FILLER_0_124_392 ();
 sg13g2_fill_2 FILLER_0_124_405 ();
 sg13g2_fill_8 FILLER_0_124_411 ();
 sg13g2_fill_8 FILLER_0_124_419 ();
 sg13g2_fill_8 FILLER_0_124_427 ();
 sg13g2_fill_1 FILLER_0_124_435 ();
 sg13g2_fill_8 FILLER_0_124_441 ();
 sg13g2_fill_8 FILLER_0_124_449 ();
 sg13g2_fill_8 FILLER_0_124_461 ();
 sg13g2_fill_8 FILLER_0_124_469 ();
 sg13g2_fill_8 FILLER_0_124_477 ();
 sg13g2_fill_8 FILLER_0_124_485 ();
 sg13g2_fill_8 FILLER_0_124_493 ();
 sg13g2_fill_8 FILLER_0_124_501 ();
 sg13g2_fill_8 FILLER_0_124_509 ();
 sg13g2_fill_4 FILLER_0_124_517 ();
 sg13g2_fill_1 FILLER_0_124_521 ();
 sg13g2_fill_2 FILLER_0_124_526 ();
 sg13g2_fill_8 FILLER_0_124_532 ();
 sg13g2_fill_2 FILLER_0_124_540 ();
 sg13g2_fill_4 FILLER_0_124_552 ();
 sg13g2_fill_4 FILLER_0_124_559 ();
 sg13g2_fill_2 FILLER_0_124_568 ();
 sg13g2_fill_2 FILLER_0_124_580 ();
 sg13g2_fill_2 FILLER_0_124_608 ();
 sg13g2_fill_1 FILLER_0_124_610 ();
 sg13g2_fill_2 FILLER_0_124_616 ();
 sg13g2_fill_2 FILLER_0_124_644 ();
 sg13g2_fill_8 FILLER_0_124_672 ();
 sg13g2_fill_8 FILLER_0_124_680 ();
 sg13g2_fill_8 FILLER_0_124_693 ();
 sg13g2_fill_8 FILLER_0_124_701 ();
 sg13g2_fill_4 FILLER_0_124_709 ();
 sg13g2_fill_2 FILLER_0_124_713 ();
 sg13g2_fill_4 FILLER_0_124_720 ();
 sg13g2_fill_2 FILLER_0_124_724 ();
 sg13g2_fill_2 FILLER_0_124_732 ();
 sg13g2_fill_1 FILLER_0_124_734 ();
 sg13g2_fill_8 FILLER_0_124_739 ();
 sg13g2_fill_4 FILLER_0_124_747 ();
 sg13g2_fill_2 FILLER_0_124_751 ();
 sg13g2_fill_1 FILLER_0_124_753 ();
 sg13g2_fill_2 FILLER_0_124_758 ();
 sg13g2_fill_1 FILLER_0_124_760 ();
 sg13g2_fill_2 FILLER_0_124_771 ();
 sg13g2_fill_4 FILLER_0_124_778 ();
 sg13g2_fill_8 FILLER_0_124_786 ();
 sg13g2_fill_8 FILLER_0_124_794 ();
 sg13g2_fill_4 FILLER_0_124_802 ();
 sg13g2_fill_2 FILLER_0_124_806 ();
 sg13g2_fill_8 FILLER_0_124_813 ();
 sg13g2_fill_8 FILLER_0_124_821 ();
 sg13g2_fill_8 FILLER_0_124_829 ();
 sg13g2_fill_2 FILLER_0_124_837 ();
 sg13g2_fill_1 FILLER_0_124_839 ();
 sg13g2_fill_2 FILLER_0_124_846 ();
 sg13g2_fill_8 FILLER_0_124_853 ();
 sg13g2_fill_4 FILLER_0_124_861 ();
 sg13g2_fill_2 FILLER_0_124_870 ();
 sg13g2_fill_2 FILLER_0_124_876 ();
 sg13g2_fill_1 FILLER_0_124_878 ();
 sg13g2_fill_2 FILLER_0_124_884 ();
 sg13g2_fill_8 FILLER_0_124_890 ();
 sg13g2_fill_4 FILLER_0_124_902 ();
 sg13g2_fill_2 FILLER_0_124_906 ();
 sg13g2_fill_8 FILLER_0_124_913 ();
 sg13g2_fill_8 FILLER_0_124_921 ();
 sg13g2_fill_2 FILLER_0_124_933 ();
 sg13g2_fill_1 FILLER_0_124_935 ();
 sg13g2_fill_8 FILLER_0_124_962 ();
 sg13g2_fill_4 FILLER_0_124_970 ();
 sg13g2_fill_1 FILLER_0_124_974 ();
 sg13g2_fill_2 FILLER_0_124_980 ();
 sg13g2_fill_4 FILLER_0_124_987 ();
 sg13g2_fill_2 FILLER_0_124_995 ();
 sg13g2_fill_1 FILLER_0_124_997 ();
 sg13g2_fill_2 FILLER_0_124_1003 ();
 sg13g2_fill_4 FILLER_0_124_1010 ();
 sg13g2_fill_8 FILLER_0_124_1017 ();
 sg13g2_fill_8 FILLER_0_124_1025 ();
 sg13g2_fill_4 FILLER_0_124_1033 ();
 sg13g2_fill_4 FILLER_0_124_1041 ();
 sg13g2_fill_4 FILLER_0_124_1050 ();
 sg13g2_fill_1 FILLER_0_124_1054 ();
 sg13g2_fill_4 FILLER_0_124_1063 ();
 sg13g2_fill_1 FILLER_0_124_1067 ();
 sg13g2_fill_4 FILLER_0_124_1075 ();
 sg13g2_fill_8 FILLER_0_124_1087 ();
 sg13g2_fill_8 FILLER_0_124_1095 ();
 sg13g2_fill_8 FILLER_0_124_1103 ();
 sg13g2_fill_4 FILLER_0_124_1111 ();
 sg13g2_fill_2 FILLER_0_124_1119 ();
 sg13g2_fill_2 FILLER_0_124_1129 ();
 sg13g2_fill_1 FILLER_0_124_1131 ();
 sg13g2_fill_2 FILLER_0_124_1137 ();
 sg13g2_fill_4 FILLER_0_124_1147 ();
 sg13g2_fill_1 FILLER_0_124_1151 ();
 sg13g2_fill_8 FILLER_0_124_1178 ();
 sg13g2_fill_4 FILLER_0_124_1186 ();
 sg13g2_fill_2 FILLER_0_124_1194 ();
 sg13g2_fill_1 FILLER_0_124_1196 ();
 sg13g2_fill_4 FILLER_0_124_1201 ();
 sg13g2_fill_2 FILLER_0_124_1210 ();
 sg13g2_fill_1 FILLER_0_124_1212 ();
 sg13g2_fill_4 FILLER_0_124_1221 ();
 sg13g2_fill_4 FILLER_0_124_1233 ();
 sg13g2_fill_2 FILLER_0_124_1237 ();
 sg13g2_fill_2 FILLER_0_124_1249 ();
 sg13g2_fill_8 FILLER_0_124_1261 ();
 sg13g2_fill_2 FILLER_0_124_1295 ();
 sg13g2_fill_8 FILLER_0_125_0 ();
 sg13g2_fill_8 FILLER_0_125_8 ();
 sg13g2_fill_8 FILLER_0_125_16 ();
 sg13g2_fill_8 FILLER_0_125_24 ();
 sg13g2_fill_8 FILLER_0_125_32 ();
 sg13g2_fill_8 FILLER_0_125_40 ();
 sg13g2_fill_8 FILLER_0_125_48 ();
 sg13g2_fill_8 FILLER_0_125_56 ();
 sg13g2_fill_8 FILLER_0_125_64 ();
 sg13g2_fill_8 FILLER_0_125_72 ();
 sg13g2_fill_8 FILLER_0_125_80 ();
 sg13g2_fill_8 FILLER_0_125_88 ();
 sg13g2_fill_8 FILLER_0_125_96 ();
 sg13g2_fill_8 FILLER_0_125_104 ();
 sg13g2_fill_8 FILLER_0_125_112 ();
 sg13g2_fill_8 FILLER_0_125_120 ();
 sg13g2_fill_8 FILLER_0_125_128 ();
 sg13g2_fill_8 FILLER_0_125_136 ();
 sg13g2_fill_8 FILLER_0_125_144 ();
 sg13g2_fill_8 FILLER_0_125_152 ();
 sg13g2_fill_8 FILLER_0_125_160 ();
 sg13g2_fill_8 FILLER_0_125_168 ();
 sg13g2_fill_8 FILLER_0_125_176 ();
 sg13g2_fill_8 FILLER_0_125_184 ();
 sg13g2_fill_8 FILLER_0_125_192 ();
 sg13g2_fill_8 FILLER_0_125_200 ();
 sg13g2_fill_8 FILLER_0_125_208 ();
 sg13g2_fill_2 FILLER_0_125_216 ();
 sg13g2_fill_1 FILLER_0_125_218 ();
 sg13g2_fill_2 FILLER_0_125_224 ();
 sg13g2_fill_8 FILLER_0_125_230 ();
 sg13g2_fill_2 FILLER_0_125_238 ();
 sg13g2_fill_1 FILLER_0_125_240 ();
 sg13g2_fill_2 FILLER_0_125_247 ();
 sg13g2_fill_8 FILLER_0_125_275 ();
 sg13g2_fill_1 FILLER_0_125_283 ();
 sg13g2_fill_8 FILLER_0_125_305 ();
 sg13g2_fill_8 FILLER_0_125_316 ();
 sg13g2_fill_4 FILLER_0_125_330 ();
 sg13g2_fill_2 FILLER_0_125_338 ();
 sg13g2_fill_8 FILLER_0_125_366 ();
 sg13g2_fill_1 FILLER_0_125_374 ();
 sg13g2_fill_2 FILLER_0_125_380 ();
 sg13g2_fill_1 FILLER_0_125_382 ();
 sg13g2_fill_8 FILLER_0_125_387 ();
 sg13g2_fill_8 FILLER_0_125_395 ();
 sg13g2_fill_8 FILLER_0_125_403 ();
 sg13g2_fill_8 FILLER_0_125_411 ();
 sg13g2_fill_8 FILLER_0_125_419 ();
 sg13g2_fill_4 FILLER_0_125_427 ();
 sg13g2_fill_1 FILLER_0_125_431 ();
 sg13g2_fill_2 FILLER_0_125_438 ();
 sg13g2_fill_8 FILLER_0_125_446 ();
 sg13g2_fill_8 FILLER_0_125_454 ();
 sg13g2_fill_8 FILLER_0_125_462 ();
 sg13g2_fill_8 FILLER_0_125_496 ();
 sg13g2_fill_4 FILLER_0_125_504 ();
 sg13g2_fill_2 FILLER_0_125_508 ();
 sg13g2_fill_1 FILLER_0_125_510 ();
 sg13g2_fill_2 FILLER_0_125_516 ();
 sg13g2_fill_8 FILLER_0_125_544 ();
 sg13g2_fill_8 FILLER_0_125_552 ();
 sg13g2_fill_4 FILLER_0_125_560 ();
 sg13g2_fill_2 FILLER_0_125_564 ();
 sg13g2_fill_1 FILLER_0_125_566 ();
 sg13g2_fill_8 FILLER_0_125_571 ();
 sg13g2_fill_1 FILLER_0_125_579 ();
 sg13g2_fill_2 FILLER_0_125_585 ();
 sg13g2_fill_8 FILLER_0_125_591 ();
 sg13g2_fill_8 FILLER_0_125_599 ();
 sg13g2_fill_8 FILLER_0_125_607 ();
 sg13g2_fill_8 FILLER_0_125_615 ();
 sg13g2_fill_2 FILLER_0_125_623 ();
 sg13g2_fill_2 FILLER_0_125_630 ();
 sg13g2_fill_1 FILLER_0_125_632 ();
 sg13g2_fill_2 FILLER_0_125_643 ();
 sg13g2_fill_2 FILLER_0_125_650 ();
 sg13g2_fill_1 FILLER_0_125_652 ();
 sg13g2_fill_4 FILLER_0_125_658 ();
 sg13g2_fill_2 FILLER_0_125_662 ();
 sg13g2_fill_1 FILLER_0_125_664 ();
 sg13g2_fill_2 FILLER_0_125_670 ();
 sg13g2_fill_8 FILLER_0_125_676 ();
 sg13g2_fill_8 FILLER_0_125_684 ();
 sg13g2_fill_8 FILLER_0_125_692 ();
 sg13g2_fill_8 FILLER_0_125_700 ();
 sg13g2_fill_8 FILLER_0_125_708 ();
 sg13g2_fill_4 FILLER_0_125_716 ();
 sg13g2_fill_8 FILLER_0_125_725 ();
 sg13g2_fill_8 FILLER_0_125_733 ();
 sg13g2_fill_4 FILLER_0_125_741 ();
 sg13g2_fill_2 FILLER_0_125_745 ();
 sg13g2_fill_2 FILLER_0_125_773 ();
 sg13g2_fill_2 FILLER_0_125_780 ();
 sg13g2_fill_8 FILLER_0_125_786 ();
 sg13g2_fill_4 FILLER_0_125_794 ();
 sg13g2_fill_2 FILLER_0_125_803 ();
 sg13g2_fill_1 FILLER_0_125_805 ();
 sg13g2_fill_2 FILLER_0_125_812 ();
 sg13g2_fill_8 FILLER_0_125_818 ();
 sg13g2_fill_8 FILLER_0_125_826 ();
 sg13g2_fill_8 FILLER_0_125_834 ();
 sg13g2_fill_8 FILLER_0_125_842 ();
 sg13g2_fill_8 FILLER_0_125_850 ();
 sg13g2_fill_8 FILLER_0_125_858 ();
 sg13g2_fill_8 FILLER_0_125_866 ();
 sg13g2_fill_4 FILLER_0_125_874 ();
 sg13g2_fill_2 FILLER_0_125_878 ();
 sg13g2_fill_1 FILLER_0_125_880 ();
 sg13g2_fill_8 FILLER_0_125_886 ();
 sg13g2_fill_8 FILLER_0_125_894 ();
 sg13g2_fill_1 FILLER_0_125_902 ();
 sg13g2_fill_8 FILLER_0_125_909 ();
 sg13g2_fill_8 FILLER_0_125_917 ();
 sg13g2_fill_4 FILLER_0_125_925 ();
 sg13g2_fill_2 FILLER_0_125_934 ();
 sg13g2_fill_2 FILLER_0_125_941 ();
 sg13g2_fill_8 FILLER_0_125_947 ();
 sg13g2_fill_2 FILLER_0_125_955 ();
 sg13g2_fill_8 FILLER_0_125_962 ();
 sg13g2_fill_8 FILLER_0_125_970 ();
 sg13g2_fill_8 FILLER_0_125_978 ();
 sg13g2_fill_8 FILLER_0_125_986 ();
 sg13g2_fill_4 FILLER_0_125_994 ();
 sg13g2_fill_2 FILLER_0_125_998 ();
 sg13g2_fill_2 FILLER_0_125_1007 ();
 sg13g2_fill_2 FILLER_0_125_1014 ();
 sg13g2_fill_8 FILLER_0_125_1020 ();
 sg13g2_fill_8 FILLER_0_125_1028 ();
 sg13g2_fill_8 FILLER_0_125_1036 ();
 sg13g2_fill_8 FILLER_0_125_1044 ();
 sg13g2_fill_8 FILLER_0_125_1052 ();
 sg13g2_fill_8 FILLER_0_125_1060 ();
 sg13g2_fill_8 FILLER_0_125_1068 ();
 sg13g2_fill_2 FILLER_0_125_1076 ();
 sg13g2_fill_1 FILLER_0_125_1078 ();
 sg13g2_fill_2 FILLER_0_125_1084 ();
 sg13g2_fill_8 FILLER_0_125_1091 ();
 sg13g2_fill_8 FILLER_0_125_1099 ();
 sg13g2_fill_8 FILLER_0_125_1107 ();
 sg13g2_fill_8 FILLER_0_125_1115 ();
 sg13g2_fill_8 FILLER_0_125_1123 ();
 sg13g2_fill_8 FILLER_0_125_1131 ();
 sg13g2_fill_4 FILLER_0_125_1139 ();
 sg13g2_fill_2 FILLER_0_125_1143 ();
 sg13g2_fill_8 FILLER_0_125_1153 ();
 sg13g2_fill_8 FILLER_0_125_1161 ();
 sg13g2_fill_1 FILLER_0_125_1169 ();
 sg13g2_fill_4 FILLER_0_125_1180 ();
 sg13g2_fill_1 FILLER_0_125_1184 ();
 sg13g2_fill_2 FILLER_0_125_1190 ();
 sg13g2_fill_4 FILLER_0_125_1200 ();
 sg13g2_fill_2 FILLER_0_125_1204 ();
 sg13g2_fill_1 FILLER_0_125_1206 ();
 sg13g2_fill_8 FILLER_0_125_1212 ();
 sg13g2_fill_4 FILLER_0_125_1220 ();
 sg13g2_fill_2 FILLER_0_125_1234 ();
 sg13g2_fill_4 FILLER_0_125_1246 ();
 sg13g2_fill_1 FILLER_0_125_1250 ();
 sg13g2_fill_2 FILLER_0_125_1277 ();
 sg13g2_fill_8 FILLER_0_125_1283 ();
 sg13g2_fill_4 FILLER_0_125_1291 ();
 sg13g2_fill_2 FILLER_0_125_1295 ();
 sg13g2_fill_8 FILLER_0_126_0 ();
 sg13g2_fill_8 FILLER_0_126_8 ();
 sg13g2_fill_8 FILLER_0_126_16 ();
 sg13g2_fill_8 FILLER_0_126_24 ();
 sg13g2_fill_8 FILLER_0_126_32 ();
 sg13g2_fill_8 FILLER_0_126_40 ();
 sg13g2_fill_8 FILLER_0_126_48 ();
 sg13g2_fill_8 FILLER_0_126_56 ();
 sg13g2_fill_8 FILLER_0_126_64 ();
 sg13g2_fill_8 FILLER_0_126_72 ();
 sg13g2_fill_8 FILLER_0_126_80 ();
 sg13g2_fill_8 FILLER_0_126_88 ();
 sg13g2_fill_8 FILLER_0_126_96 ();
 sg13g2_fill_8 FILLER_0_126_104 ();
 sg13g2_fill_8 FILLER_0_126_112 ();
 sg13g2_fill_8 FILLER_0_126_120 ();
 sg13g2_fill_8 FILLER_0_126_128 ();
 sg13g2_fill_8 FILLER_0_126_136 ();
 sg13g2_fill_8 FILLER_0_126_144 ();
 sg13g2_fill_8 FILLER_0_126_152 ();
 sg13g2_fill_8 FILLER_0_126_160 ();
 sg13g2_fill_8 FILLER_0_126_168 ();
 sg13g2_fill_8 FILLER_0_126_176 ();
 sg13g2_fill_8 FILLER_0_126_184 ();
 sg13g2_fill_8 FILLER_0_126_192 ();
 sg13g2_fill_4 FILLER_0_126_200 ();
 sg13g2_fill_2 FILLER_0_126_204 ();
 sg13g2_fill_1 FILLER_0_126_206 ();
 sg13g2_fill_8 FILLER_0_126_233 ();
 sg13g2_fill_1 FILLER_0_126_241 ();
 sg13g2_fill_2 FILLER_0_126_247 ();
 sg13g2_fill_4 FILLER_0_126_270 ();
 sg13g2_fill_2 FILLER_0_126_274 ();
 sg13g2_fill_8 FILLER_0_126_302 ();
 sg13g2_fill_8 FILLER_0_126_310 ();
 sg13g2_fill_2 FILLER_0_126_318 ();
 sg13g2_fill_1 FILLER_0_126_320 ();
 sg13g2_fill_8 FILLER_0_126_347 ();
 sg13g2_fill_4 FILLER_0_126_355 ();
 sg13g2_fill_2 FILLER_0_126_359 ();
 sg13g2_fill_8 FILLER_0_126_382 ();
 sg13g2_fill_4 FILLER_0_126_390 ();
 sg13g2_fill_1 FILLER_0_126_394 ();
 sg13g2_fill_4 FILLER_0_126_400 ();
 sg13g2_fill_1 FILLER_0_126_404 ();
 sg13g2_fill_2 FILLER_0_126_409 ();
 sg13g2_fill_2 FILLER_0_126_416 ();
 sg13g2_fill_4 FILLER_0_126_422 ();
 sg13g2_fill_2 FILLER_0_126_431 ();
 sg13g2_fill_2 FILLER_0_126_437 ();
 sg13g2_fill_8 FILLER_0_126_445 ();
 sg13g2_fill_8 FILLER_0_126_453 ();
 sg13g2_fill_8 FILLER_0_126_461 ();
 sg13g2_fill_8 FILLER_0_126_469 ();
 sg13g2_fill_4 FILLER_0_126_477 ();
 sg13g2_fill_8 FILLER_0_126_507 ();
 sg13g2_fill_8 FILLER_0_126_515 ();
 sg13g2_fill_1 FILLER_0_126_523 ();
 sg13g2_fill_8 FILLER_0_126_529 ();
 sg13g2_fill_8 FILLER_0_126_537 ();
 sg13g2_fill_8 FILLER_0_126_545 ();
 sg13g2_fill_8 FILLER_0_126_553 ();
 sg13g2_fill_8 FILLER_0_126_561 ();
 sg13g2_fill_8 FILLER_0_126_569 ();
 sg13g2_fill_8 FILLER_0_126_577 ();
 sg13g2_fill_8 FILLER_0_126_585 ();
 sg13g2_fill_8 FILLER_0_126_593 ();
 sg13g2_fill_8 FILLER_0_126_601 ();
 sg13g2_fill_8 FILLER_0_126_609 ();
 sg13g2_fill_8 FILLER_0_126_617 ();
 sg13g2_fill_1 FILLER_0_126_625 ();
 sg13g2_fill_2 FILLER_0_126_632 ();
 sg13g2_fill_4 FILLER_0_126_639 ();
 sg13g2_fill_2 FILLER_0_126_643 ();
 sg13g2_fill_1 FILLER_0_126_645 ();
 sg13g2_fill_2 FILLER_0_126_672 ();
 sg13g2_fill_8 FILLER_0_126_680 ();
 sg13g2_fill_8 FILLER_0_126_688 ();
 sg13g2_fill_8 FILLER_0_126_696 ();
 sg13g2_fill_8 FILLER_0_126_704 ();
 sg13g2_fill_4 FILLER_0_126_712 ();
 sg13g2_fill_2 FILLER_0_126_716 ();
 sg13g2_fill_1 FILLER_0_126_718 ();
 sg13g2_fill_2 FILLER_0_126_724 ();
 sg13g2_fill_8 FILLER_0_126_730 ();
 sg13g2_fill_4 FILLER_0_126_738 ();
 sg13g2_fill_2 FILLER_0_126_742 ();
 sg13g2_fill_1 FILLER_0_126_744 ();
 sg13g2_fill_2 FILLER_0_126_750 ();
 sg13g2_fill_8 FILLER_0_126_757 ();
 sg13g2_fill_8 FILLER_0_126_765 ();
 sg13g2_fill_8 FILLER_0_126_773 ();
 sg13g2_fill_8 FILLER_0_126_781 ();
 sg13g2_fill_2 FILLER_0_126_789 ();
 sg13g2_fill_2 FILLER_0_126_817 ();
 sg13g2_fill_8 FILLER_0_126_825 ();
 sg13g2_fill_8 FILLER_0_126_833 ();
 sg13g2_fill_2 FILLER_0_126_841 ();
 sg13g2_fill_8 FILLER_0_126_869 ();
 sg13g2_fill_1 FILLER_0_126_877 ();
 sg13g2_fill_8 FILLER_0_126_884 ();
 sg13g2_fill_4 FILLER_0_126_902 ();
 sg13g2_fill_8 FILLER_0_126_912 ();
 sg13g2_fill_8 FILLER_0_126_920 ();
 sg13g2_fill_4 FILLER_0_126_928 ();
 sg13g2_fill_2 FILLER_0_126_932 ();
 sg13g2_fill_1 FILLER_0_126_934 ();
 sg13g2_fill_2 FILLER_0_126_961 ();
 sg13g2_fill_8 FILLER_0_126_969 ();
 sg13g2_fill_8 FILLER_0_126_977 ();
 sg13g2_fill_1 FILLER_0_126_985 ();
 sg13g2_fill_8 FILLER_0_126_991 ();
 sg13g2_fill_8 FILLER_0_126_999 ();
 sg13g2_fill_8 FILLER_0_126_1007 ();
 sg13g2_fill_8 FILLER_0_126_1015 ();
 sg13g2_fill_8 FILLER_0_126_1023 ();
 sg13g2_fill_8 FILLER_0_126_1035 ();
 sg13g2_fill_8 FILLER_0_126_1043 ();
 sg13g2_fill_8 FILLER_0_126_1051 ();
 sg13g2_fill_8 FILLER_0_126_1059 ();
 sg13g2_fill_8 FILLER_0_126_1067 ();
 sg13g2_fill_2 FILLER_0_126_1075 ();
 sg13g2_fill_1 FILLER_0_126_1077 ();
 sg13g2_fill_8 FILLER_0_126_1084 ();
 sg13g2_fill_8 FILLER_0_126_1092 ();
 sg13g2_fill_8 FILLER_0_126_1100 ();
 sg13g2_fill_8 FILLER_0_126_1108 ();
 sg13g2_fill_4 FILLER_0_126_1116 ();
 sg13g2_fill_1 FILLER_0_126_1120 ();
 sg13g2_fill_8 FILLER_0_126_1147 ();
 sg13g2_fill_8 FILLER_0_126_1155 ();
 sg13g2_fill_8 FILLER_0_126_1163 ();
 sg13g2_fill_2 FILLER_0_126_1171 ();
 sg13g2_fill_2 FILLER_0_126_1177 ();
 sg13g2_fill_2 FILLER_0_126_1205 ();
 sg13g2_fill_2 FILLER_0_126_1213 ();
 sg13g2_fill_8 FILLER_0_126_1220 ();
 sg13g2_fill_2 FILLER_0_126_1228 ();
 sg13g2_fill_1 FILLER_0_126_1230 ();
 sg13g2_fill_8 FILLER_0_126_1236 ();
 sg13g2_fill_8 FILLER_0_126_1244 ();
 sg13g2_fill_8 FILLER_0_126_1252 ();
 sg13g2_fill_8 FILLER_0_126_1260 ();
 sg13g2_fill_8 FILLER_0_126_1268 ();
 sg13g2_fill_8 FILLER_0_126_1284 ();
 sg13g2_fill_4 FILLER_0_126_1292 ();
 sg13g2_fill_1 FILLER_0_126_1296 ();
 sg13g2_fill_8 FILLER_0_127_0 ();
 sg13g2_fill_8 FILLER_0_127_8 ();
 sg13g2_fill_8 FILLER_0_127_16 ();
 sg13g2_fill_8 FILLER_0_127_24 ();
 sg13g2_fill_8 FILLER_0_127_32 ();
 sg13g2_fill_8 FILLER_0_127_40 ();
 sg13g2_fill_8 FILLER_0_127_48 ();
 sg13g2_fill_8 FILLER_0_127_56 ();
 sg13g2_fill_8 FILLER_0_127_64 ();
 sg13g2_fill_8 FILLER_0_127_72 ();
 sg13g2_fill_8 FILLER_0_127_80 ();
 sg13g2_fill_8 FILLER_0_127_88 ();
 sg13g2_fill_8 FILLER_0_127_96 ();
 sg13g2_fill_8 FILLER_0_127_104 ();
 sg13g2_fill_8 FILLER_0_127_112 ();
 sg13g2_fill_8 FILLER_0_127_120 ();
 sg13g2_fill_8 FILLER_0_127_128 ();
 sg13g2_fill_8 FILLER_0_127_136 ();
 sg13g2_fill_8 FILLER_0_127_144 ();
 sg13g2_fill_8 FILLER_0_127_152 ();
 sg13g2_fill_8 FILLER_0_127_160 ();
 sg13g2_fill_8 FILLER_0_127_168 ();
 sg13g2_fill_8 FILLER_0_127_176 ();
 sg13g2_fill_8 FILLER_0_127_184 ();
 sg13g2_fill_8 FILLER_0_127_192 ();
 sg13g2_fill_8 FILLER_0_127_200 ();
 sg13g2_fill_8 FILLER_0_127_208 ();
 sg13g2_fill_8 FILLER_0_127_216 ();
 sg13g2_fill_8 FILLER_0_127_224 ();
 sg13g2_fill_1 FILLER_0_127_232 ();
 sg13g2_fill_2 FILLER_0_127_238 ();
 sg13g2_fill_1 FILLER_0_127_240 ();
 sg13g2_fill_2 FILLER_0_127_245 ();
 sg13g2_fill_2 FILLER_0_127_252 ();
 sg13g2_fill_8 FILLER_0_127_258 ();
 sg13g2_fill_8 FILLER_0_127_266 ();
 sg13g2_fill_2 FILLER_0_127_274 ();
 sg13g2_fill_1 FILLER_0_127_276 ();
 sg13g2_fill_2 FILLER_0_127_281 ();
 sg13g2_fill_8 FILLER_0_127_288 ();
 sg13g2_fill_8 FILLER_0_127_296 ();
 sg13g2_fill_8 FILLER_0_127_304 ();
 sg13g2_fill_4 FILLER_0_127_312 ();
 sg13g2_fill_1 FILLER_0_127_316 ();
 sg13g2_fill_8 FILLER_0_127_322 ();
 sg13g2_fill_4 FILLER_0_127_334 ();
 sg13g2_fill_2 FILLER_0_127_338 ();
 sg13g2_fill_1 FILLER_0_127_340 ();
 sg13g2_fill_8 FILLER_0_127_346 ();
 sg13g2_fill_8 FILLER_0_127_354 ();
 sg13g2_fill_2 FILLER_0_127_362 ();
 sg13g2_fill_1 FILLER_0_127_364 ();
 sg13g2_fill_8 FILLER_0_127_370 ();
 sg13g2_fill_8 FILLER_0_127_378 ();
 sg13g2_fill_4 FILLER_0_127_386 ();
 sg13g2_fill_2 FILLER_0_127_390 ();
 sg13g2_fill_1 FILLER_0_127_392 ();
 sg13g2_fill_8 FILLER_0_127_398 ();
 sg13g2_fill_2 FILLER_0_127_406 ();
 sg13g2_fill_1 FILLER_0_127_408 ();
 sg13g2_fill_8 FILLER_0_127_435 ();
 sg13g2_fill_8 FILLER_0_127_443 ();
 sg13g2_fill_8 FILLER_0_127_451 ();
 sg13g2_fill_4 FILLER_0_127_459 ();
 sg13g2_fill_2 FILLER_0_127_463 ();
 sg13g2_fill_1 FILLER_0_127_465 ();
 sg13g2_fill_2 FILLER_0_127_471 ();
 sg13g2_fill_2 FILLER_0_127_477 ();
 sg13g2_fill_8 FILLER_0_127_484 ();
 sg13g2_fill_1 FILLER_0_127_492 ();
 sg13g2_fill_2 FILLER_0_127_497 ();
 sg13g2_fill_8 FILLER_0_127_504 ();
 sg13g2_fill_8 FILLER_0_127_512 ();
 sg13g2_fill_4 FILLER_0_127_520 ();
 sg13g2_fill_2 FILLER_0_127_524 ();
 sg13g2_fill_1 FILLER_0_127_526 ();
 sg13g2_fill_8 FILLER_0_127_553 ();
 sg13g2_fill_8 FILLER_0_127_561 ();
 sg13g2_fill_8 FILLER_0_127_569 ();
 sg13g2_fill_4 FILLER_0_127_577 ();
 sg13g2_fill_2 FILLER_0_127_581 ();
 sg13g2_fill_1 FILLER_0_127_583 ();
 sg13g2_fill_8 FILLER_0_127_589 ();
 sg13g2_fill_8 FILLER_0_127_597 ();
 sg13g2_fill_4 FILLER_0_127_605 ();
 sg13g2_fill_1 FILLER_0_127_609 ();
 sg13g2_fill_8 FILLER_0_127_615 ();
 sg13g2_fill_8 FILLER_0_127_623 ();
 sg13g2_fill_8 FILLER_0_127_631 ();
 sg13g2_fill_4 FILLER_0_127_639 ();
 sg13g2_fill_1 FILLER_0_127_643 ();
 sg13g2_fill_2 FILLER_0_127_670 ();
 sg13g2_fill_8 FILLER_0_127_677 ();
 sg13g2_fill_2 FILLER_0_127_685 ();
 sg13g2_fill_1 FILLER_0_127_687 ();
 sg13g2_fill_4 FILLER_0_127_693 ();
 sg13g2_fill_1 FILLER_0_127_697 ();
 sg13g2_fill_8 FILLER_0_127_702 ();
 sg13g2_fill_4 FILLER_0_127_710 ();
 sg13g2_fill_2 FILLER_0_127_714 ();
 sg13g2_fill_2 FILLER_0_127_742 ();
 sg13g2_fill_2 FILLER_0_127_749 ();
 sg13g2_fill_1 FILLER_0_127_751 ();
 sg13g2_fill_8 FILLER_0_127_758 ();
 sg13g2_fill_8 FILLER_0_127_766 ();
 sg13g2_fill_4 FILLER_0_127_774 ();
 sg13g2_fill_8 FILLER_0_127_783 ();
 sg13g2_fill_8 FILLER_0_127_791 ();
 sg13g2_fill_2 FILLER_0_127_799 ();
 sg13g2_fill_4 FILLER_0_127_805 ();
 sg13g2_fill_1 FILLER_0_127_809 ();
 sg13g2_fill_2 FILLER_0_127_815 ();
 sg13g2_fill_8 FILLER_0_127_822 ();
 sg13g2_fill_8 FILLER_0_127_830 ();
 sg13g2_fill_8 FILLER_0_127_838 ();
 sg13g2_fill_4 FILLER_0_127_846 ();
 sg13g2_fill_2 FILLER_0_127_850 ();
 sg13g2_fill_2 FILLER_0_127_857 ();
 sg13g2_fill_8 FILLER_0_127_866 ();
 sg13g2_fill_2 FILLER_0_127_874 ();
 sg13g2_fill_4 FILLER_0_127_881 ();
 sg13g2_fill_2 FILLER_0_127_885 ();
 sg13g2_fill_1 FILLER_0_127_887 ();
 sg13g2_fill_8 FILLER_0_127_892 ();
 sg13g2_fill_1 FILLER_0_127_900 ();
 sg13g2_fill_8 FILLER_0_127_909 ();
 sg13g2_fill_8 FILLER_0_127_917 ();
 sg13g2_fill_4 FILLER_0_127_925 ();
 sg13g2_fill_2 FILLER_0_127_929 ();
 sg13g2_fill_1 FILLER_0_127_931 ();
 sg13g2_fill_8 FILLER_0_127_937 ();
 sg13g2_fill_4 FILLER_0_127_945 ();
 sg13g2_fill_8 FILLER_0_127_954 ();
 sg13g2_fill_8 FILLER_0_127_962 ();
 sg13g2_fill_4 FILLER_0_127_970 ();
 sg13g2_fill_2 FILLER_0_127_974 ();
 sg13g2_fill_8 FILLER_0_127_981 ();
 sg13g2_fill_8 FILLER_0_127_989 ();
 sg13g2_fill_8 FILLER_0_127_997 ();
 sg13g2_fill_4 FILLER_0_127_1005 ();
 sg13g2_fill_2 FILLER_0_127_1015 ();
 sg13g2_fill_8 FILLER_0_127_1026 ();
 sg13g2_fill_4 FILLER_0_127_1034 ();
 sg13g2_fill_2 FILLER_0_127_1038 ();
 sg13g2_fill_2 FILLER_0_127_1044 ();
 sg13g2_fill_2 FILLER_0_127_1051 ();
 sg13g2_fill_2 FILLER_0_127_1057 ();
 sg13g2_fill_2 FILLER_0_127_1065 ();
 sg13g2_fill_1 FILLER_0_127_1067 ();
 sg13g2_fill_2 FILLER_0_127_1072 ();
 sg13g2_fill_1 FILLER_0_127_1074 ();
 sg13g2_fill_2 FILLER_0_127_1080 ();
 sg13g2_fill_1 FILLER_0_127_1082 ();
 sg13g2_fill_2 FILLER_0_127_1089 ();
 sg13g2_fill_8 FILLER_0_127_1095 ();
 sg13g2_fill_8 FILLER_0_127_1103 ();
 sg13g2_fill_2 FILLER_0_127_1111 ();
 sg13g2_fill_2 FILLER_0_127_1123 ();
 sg13g2_fill_4 FILLER_0_127_1135 ();
 sg13g2_fill_1 FILLER_0_127_1139 ();
 sg13g2_fill_4 FILLER_0_127_1145 ();
 sg13g2_fill_2 FILLER_0_127_1155 ();
 sg13g2_fill_2 FILLER_0_127_1162 ();
 sg13g2_fill_8 FILLER_0_127_1169 ();
 sg13g2_fill_8 FILLER_0_127_1177 ();
 sg13g2_fill_4 FILLER_0_127_1185 ();
 sg13g2_fill_2 FILLER_0_127_1194 ();
 sg13g2_fill_8 FILLER_0_127_1201 ();
 sg13g2_fill_8 FILLER_0_127_1209 ();
 sg13g2_fill_4 FILLER_0_127_1217 ();
 sg13g2_fill_1 FILLER_0_127_1221 ();
 sg13g2_fill_8 FILLER_0_127_1230 ();
 sg13g2_fill_8 FILLER_0_127_1238 ();
 sg13g2_fill_8 FILLER_0_127_1246 ();
 sg13g2_fill_8 FILLER_0_127_1254 ();
 sg13g2_fill_8 FILLER_0_127_1262 ();
 sg13g2_fill_8 FILLER_0_127_1270 ();
 sg13g2_fill_8 FILLER_0_127_1278 ();
 sg13g2_fill_8 FILLER_0_127_1286 ();
 sg13g2_fill_2 FILLER_0_127_1294 ();
 sg13g2_fill_1 FILLER_0_127_1296 ();
 sg13g2_fill_8 FILLER_0_128_0 ();
 sg13g2_fill_8 FILLER_0_128_8 ();
 sg13g2_fill_8 FILLER_0_128_16 ();
 sg13g2_fill_8 FILLER_0_128_24 ();
 sg13g2_fill_8 FILLER_0_128_32 ();
 sg13g2_fill_8 FILLER_0_128_40 ();
 sg13g2_fill_8 FILLER_0_128_48 ();
 sg13g2_fill_8 FILLER_0_128_56 ();
 sg13g2_fill_8 FILLER_0_128_64 ();
 sg13g2_fill_8 FILLER_0_128_72 ();
 sg13g2_fill_8 FILLER_0_128_80 ();
 sg13g2_fill_8 FILLER_0_128_88 ();
 sg13g2_fill_8 FILLER_0_128_96 ();
 sg13g2_fill_8 FILLER_0_128_104 ();
 sg13g2_fill_8 FILLER_0_128_112 ();
 sg13g2_fill_8 FILLER_0_128_120 ();
 sg13g2_fill_8 FILLER_0_128_128 ();
 sg13g2_fill_8 FILLER_0_128_136 ();
 sg13g2_fill_8 FILLER_0_128_144 ();
 sg13g2_fill_8 FILLER_0_128_152 ();
 sg13g2_fill_8 FILLER_0_128_160 ();
 sg13g2_fill_8 FILLER_0_128_168 ();
 sg13g2_fill_8 FILLER_0_128_176 ();
 sg13g2_fill_8 FILLER_0_128_184 ();
 sg13g2_fill_8 FILLER_0_128_192 ();
 sg13g2_fill_8 FILLER_0_128_200 ();
 sg13g2_fill_8 FILLER_0_128_208 ();
 sg13g2_fill_4 FILLER_0_128_216 ();
 sg13g2_fill_2 FILLER_0_128_220 ();
 sg13g2_fill_8 FILLER_0_128_248 ();
 sg13g2_fill_8 FILLER_0_128_256 ();
 sg13g2_fill_8 FILLER_0_128_264 ();
 sg13g2_fill_8 FILLER_0_128_272 ();
 sg13g2_fill_8 FILLER_0_128_280 ();
 sg13g2_fill_8 FILLER_0_128_288 ();
 sg13g2_fill_4 FILLER_0_128_296 ();
 sg13g2_fill_2 FILLER_0_128_300 ();
 sg13g2_fill_8 FILLER_0_128_306 ();
 sg13g2_fill_8 FILLER_0_128_314 ();
 sg13g2_fill_8 FILLER_0_128_322 ();
 sg13g2_fill_8 FILLER_0_128_330 ();
 sg13g2_fill_1 FILLER_0_128_338 ();
 sg13g2_fill_2 FILLER_0_128_345 ();
 sg13g2_fill_8 FILLER_0_128_373 ();
 sg13g2_fill_8 FILLER_0_128_381 ();
 sg13g2_fill_4 FILLER_0_128_389 ();
 sg13g2_fill_1 FILLER_0_128_393 ();
 sg13g2_fill_2 FILLER_0_128_399 ();
 sg13g2_fill_4 FILLER_0_128_427 ();
 sg13g2_fill_1 FILLER_0_128_431 ();
 sg13g2_fill_2 FILLER_0_128_437 ();
 sg13g2_fill_8 FILLER_0_128_444 ();
 sg13g2_fill_8 FILLER_0_128_452 ();
 sg13g2_fill_8 FILLER_0_128_460 ();
 sg13g2_fill_8 FILLER_0_128_468 ();
 sg13g2_fill_2 FILLER_0_128_476 ();
 sg13g2_fill_1 FILLER_0_128_478 ();
 sg13g2_fill_8 FILLER_0_128_484 ();
 sg13g2_fill_8 FILLER_0_128_492 ();
 sg13g2_fill_8 FILLER_0_128_500 ();
 sg13g2_fill_8 FILLER_0_128_508 ();
 sg13g2_fill_8 FILLER_0_128_516 ();
 sg13g2_fill_8 FILLER_0_128_524 ();
 sg13g2_fill_4 FILLER_0_128_532 ();
 sg13g2_fill_2 FILLER_0_128_536 ();
 sg13g2_fill_8 FILLER_0_128_559 ();
 sg13g2_fill_8 FILLER_0_128_567 ();
 sg13g2_fill_2 FILLER_0_128_575 ();
 sg13g2_fill_1 FILLER_0_128_577 ();
 sg13g2_fill_2 FILLER_0_128_583 ();
 sg13g2_fill_2 FILLER_0_128_591 ();
 sg13g2_fill_2 FILLER_0_128_619 ();
 sg13g2_fill_2 FILLER_0_128_626 ();
 sg13g2_fill_2 FILLER_0_128_632 ();
 sg13g2_fill_1 FILLER_0_128_634 ();
 sg13g2_fill_2 FILLER_0_128_640 ();
 sg13g2_fill_2 FILLER_0_128_647 ();
 sg13g2_fill_8 FILLER_0_128_653 ();
 sg13g2_fill_8 FILLER_0_128_661 ();
 sg13g2_fill_8 FILLER_0_128_669 ();
 sg13g2_fill_8 FILLER_0_128_677 ();
 sg13g2_fill_4 FILLER_0_128_685 ();
 sg13g2_fill_8 FILLER_0_128_715 ();
 sg13g2_fill_8 FILLER_0_128_727 ();
 sg13g2_fill_2 FILLER_0_128_735 ();
 sg13g2_fill_1 FILLER_0_128_737 ();
 sg13g2_fill_4 FILLER_0_128_742 ();
 sg13g2_fill_4 FILLER_0_128_751 ();
 sg13g2_fill_8 FILLER_0_128_781 ();
 sg13g2_fill_4 FILLER_0_128_794 ();
 sg13g2_fill_1 FILLER_0_128_798 ();
 sg13g2_fill_2 FILLER_0_128_804 ();
 sg13g2_fill_8 FILLER_0_128_811 ();
 sg13g2_fill_8 FILLER_0_128_819 ();
 sg13g2_fill_4 FILLER_0_128_827 ();
 sg13g2_fill_2 FILLER_0_128_836 ();
 sg13g2_fill_2 FILLER_0_128_842 ();
 sg13g2_fill_1 FILLER_0_128_844 ();
 sg13g2_fill_8 FILLER_0_128_850 ();
 sg13g2_fill_8 FILLER_0_128_858 ();
 sg13g2_fill_2 FILLER_0_128_871 ();
 sg13g2_fill_2 FILLER_0_128_877 ();
 sg13g2_fill_8 FILLER_0_128_905 ();
 sg13g2_fill_4 FILLER_0_128_913 ();
 sg13g2_fill_2 FILLER_0_128_917 ();
 sg13g2_fill_8 FILLER_0_128_945 ();
 sg13g2_fill_2 FILLER_0_128_953 ();
 sg13g2_fill_1 FILLER_0_128_955 ();
 sg13g2_fill_2 FILLER_0_128_960 ();
 sg13g2_fill_8 FILLER_0_128_966 ();
 sg13g2_fill_4 FILLER_0_128_974 ();
 sg13g2_fill_1 FILLER_0_128_978 ();
 sg13g2_fill_2 FILLER_0_128_991 ();
 sg13g2_fill_2 FILLER_0_128_998 ();
 sg13g2_fill_2 FILLER_0_128_1004 ();
 sg13g2_fill_2 FILLER_0_128_1011 ();
 sg13g2_fill_2 FILLER_0_128_1025 ();
 sg13g2_fill_2 FILLER_0_128_1033 ();
 sg13g2_fill_2 FILLER_0_128_1040 ();
 sg13g2_fill_8 FILLER_0_128_1047 ();
 sg13g2_fill_4 FILLER_0_128_1055 ();
 sg13g2_fill_2 FILLER_0_128_1059 ();
 sg13g2_fill_1 FILLER_0_128_1061 ();
 sg13g2_fill_2 FILLER_0_128_1067 ();
 sg13g2_fill_2 FILLER_0_128_1074 ();
 sg13g2_fill_4 FILLER_0_128_1083 ();
 sg13g2_fill_8 FILLER_0_128_1095 ();
 sg13g2_fill_8 FILLER_0_128_1103 ();
 sg13g2_fill_8 FILLER_0_128_1111 ();
 sg13g2_fill_8 FILLER_0_128_1119 ();
 sg13g2_fill_8 FILLER_0_128_1127 ();
 sg13g2_fill_4 FILLER_0_128_1135 ();
 sg13g2_fill_2 FILLER_0_128_1139 ();
 sg13g2_fill_4 FILLER_0_128_1146 ();
 sg13g2_fill_8 FILLER_0_128_1155 ();
 sg13g2_fill_8 FILLER_0_128_1163 ();
 sg13g2_fill_8 FILLER_0_128_1171 ();
 sg13g2_fill_8 FILLER_0_128_1179 ();
 sg13g2_fill_8 FILLER_0_128_1187 ();
 sg13g2_fill_8 FILLER_0_128_1200 ();
 sg13g2_fill_8 FILLER_0_128_1208 ();
 sg13g2_fill_8 FILLER_0_128_1216 ();
 sg13g2_fill_8 FILLER_0_128_1224 ();
 sg13g2_fill_4 FILLER_0_128_1232 ();
 sg13g2_fill_2 FILLER_0_128_1236 ();
 sg13g2_fill_8 FILLER_0_128_1264 ();
 sg13g2_fill_8 FILLER_0_128_1272 ();
 sg13g2_fill_2 FILLER_0_128_1285 ();
 sg13g2_fill_4 FILLER_0_128_1291 ();
 sg13g2_fill_2 FILLER_0_128_1295 ();
 sg13g2_fill_8 FILLER_0_129_0 ();
 sg13g2_fill_8 FILLER_0_129_8 ();
 sg13g2_fill_8 FILLER_0_129_16 ();
 sg13g2_fill_8 FILLER_0_129_24 ();
 sg13g2_fill_8 FILLER_0_129_32 ();
 sg13g2_fill_8 FILLER_0_129_40 ();
 sg13g2_fill_8 FILLER_0_129_48 ();
 sg13g2_fill_8 FILLER_0_129_56 ();
 sg13g2_fill_8 FILLER_0_129_64 ();
 sg13g2_fill_8 FILLER_0_129_72 ();
 sg13g2_fill_8 FILLER_0_129_80 ();
 sg13g2_fill_8 FILLER_0_129_88 ();
 sg13g2_fill_8 FILLER_0_129_96 ();
 sg13g2_fill_8 FILLER_0_129_104 ();
 sg13g2_fill_8 FILLER_0_129_112 ();
 sg13g2_fill_8 FILLER_0_129_120 ();
 sg13g2_fill_8 FILLER_0_129_128 ();
 sg13g2_fill_8 FILLER_0_129_136 ();
 sg13g2_fill_8 FILLER_0_129_144 ();
 sg13g2_fill_8 FILLER_0_129_152 ();
 sg13g2_fill_8 FILLER_0_129_160 ();
 sg13g2_fill_8 FILLER_0_129_168 ();
 sg13g2_fill_8 FILLER_0_129_176 ();
 sg13g2_fill_8 FILLER_0_129_184 ();
 sg13g2_fill_8 FILLER_0_129_192 ();
 sg13g2_fill_8 FILLER_0_129_200 ();
 sg13g2_fill_8 FILLER_0_129_208 ();
 sg13g2_fill_8 FILLER_0_129_216 ();
 sg13g2_fill_8 FILLER_0_129_224 ();
 sg13g2_fill_8 FILLER_0_129_232 ();
 sg13g2_fill_8 FILLER_0_129_240 ();
 sg13g2_fill_8 FILLER_0_129_248 ();
 sg13g2_fill_8 FILLER_0_129_256 ();
 sg13g2_fill_8 FILLER_0_129_264 ();
 sg13g2_fill_8 FILLER_0_129_272 ();
 sg13g2_fill_8 FILLER_0_129_280 ();
 sg13g2_fill_4 FILLER_0_129_288 ();
 sg13g2_fill_2 FILLER_0_129_292 ();
 sg13g2_fill_2 FILLER_0_129_299 ();
 sg13g2_fill_4 FILLER_0_129_306 ();
 sg13g2_fill_2 FILLER_0_129_310 ();
 sg13g2_fill_2 FILLER_0_129_317 ();
 sg13g2_fill_4 FILLER_0_129_325 ();
 sg13g2_fill_1 FILLER_0_129_329 ();
 sg13g2_fill_2 FILLER_0_129_335 ();
 sg13g2_fill_2 FILLER_0_129_345 ();
 sg13g2_fill_4 FILLER_0_129_352 ();
 sg13g2_fill_2 FILLER_0_129_356 ();
 sg13g2_fill_1 FILLER_0_129_358 ();
 sg13g2_fill_2 FILLER_0_129_385 ();
 sg13g2_fill_1 FILLER_0_129_387 ();
 sg13g2_fill_2 FILLER_0_129_393 ();
 sg13g2_fill_1 FILLER_0_129_395 ();
 sg13g2_fill_8 FILLER_0_129_400 ();
 sg13g2_fill_2 FILLER_0_129_408 ();
 sg13g2_fill_1 FILLER_0_129_410 ();
 sg13g2_fill_4 FILLER_0_129_419 ();
 sg13g2_fill_2 FILLER_0_129_423 ();
 sg13g2_fill_4 FILLER_0_129_446 ();
 sg13g2_fill_2 FILLER_0_129_450 ();
 sg13g2_fill_1 FILLER_0_129_452 ();
 sg13g2_fill_8 FILLER_0_129_460 ();
 sg13g2_fill_4 FILLER_0_129_468 ();
 sg13g2_fill_2 FILLER_0_129_472 ();
 sg13g2_fill_1 FILLER_0_129_474 ();
 sg13g2_fill_8 FILLER_0_129_480 ();
 sg13g2_fill_1 FILLER_0_129_488 ();
 sg13g2_fill_8 FILLER_0_129_510 ();
 sg13g2_fill_4 FILLER_0_129_544 ();
 sg13g2_fill_4 FILLER_0_129_552 ();
 sg13g2_fill_2 FILLER_0_129_582 ();
 sg13g2_fill_2 FILLER_0_129_588 ();
 sg13g2_fill_2 FILLER_0_129_595 ();
 sg13g2_fill_8 FILLER_0_129_600 ();
 sg13g2_fill_1 FILLER_0_129_608 ();
 sg13g2_fill_4 FILLER_0_129_615 ();
 sg13g2_fill_4 FILLER_0_129_624 ();
 sg13g2_fill_2 FILLER_0_129_628 ();
 sg13g2_fill_1 FILLER_0_129_630 ();
 sg13g2_fill_8 FILLER_0_129_637 ();
 sg13g2_fill_8 FILLER_0_129_645 ();
 sg13g2_fill_8 FILLER_0_129_653 ();
 sg13g2_fill_8 FILLER_0_129_661 ();
 sg13g2_fill_4 FILLER_0_129_669 ();
 sg13g2_fill_2 FILLER_0_129_673 ();
 sg13g2_fill_8 FILLER_0_129_680 ();
 sg13g2_fill_8 FILLER_0_129_688 ();
 sg13g2_fill_8 FILLER_0_129_701 ();
 sg13g2_fill_8 FILLER_0_129_714 ();
 sg13g2_fill_2 FILLER_0_129_727 ();
 sg13g2_fill_4 FILLER_0_129_755 ();
 sg13g2_fill_2 FILLER_0_129_759 ();
 sg13g2_fill_2 FILLER_0_129_765 ();
 sg13g2_fill_2 FILLER_0_129_775 ();
 sg13g2_fill_4 FILLER_0_129_782 ();
 sg13g2_fill_2 FILLER_0_129_790 ();
 sg13g2_fill_8 FILLER_0_129_818 ();
 sg13g2_fill_4 FILLER_0_129_826 ();
 sg13g2_fill_2 FILLER_0_129_830 ();
 sg13g2_fill_8 FILLER_0_129_858 ();
 sg13g2_fill_8 FILLER_0_129_866 ();
 sg13g2_fill_2 FILLER_0_129_874 ();
 sg13g2_fill_4 FILLER_0_129_881 ();
 sg13g2_fill_2 FILLER_0_129_885 ();
 sg13g2_fill_1 FILLER_0_129_887 ();
 sg13g2_fill_2 FILLER_0_129_914 ();
 sg13g2_fill_8 FILLER_0_129_937 ();
 sg13g2_fill_8 FILLER_0_129_945 ();
 sg13g2_fill_1 FILLER_0_129_953 ();
 sg13g2_fill_2 FILLER_0_129_958 ();
 sg13g2_fill_8 FILLER_0_129_965 ();
 sg13g2_fill_8 FILLER_0_129_973 ();
 sg13g2_fill_8 FILLER_0_129_981 ();
 sg13g2_fill_8 FILLER_0_129_989 ();
 sg13g2_fill_8 FILLER_0_129_997 ();
 sg13g2_fill_8 FILLER_0_129_1005 ();
 sg13g2_fill_8 FILLER_0_129_1013 ();
 sg13g2_fill_8 FILLER_0_129_1021 ();
 sg13g2_fill_8 FILLER_0_129_1029 ();
 sg13g2_fill_8 FILLER_0_129_1037 ();
 sg13g2_fill_8 FILLER_0_129_1045 ();
 sg13g2_fill_2 FILLER_0_129_1053 ();
 sg13g2_fill_2 FILLER_0_129_1061 ();
 sg13g2_fill_2 FILLER_0_129_1068 ();
 sg13g2_fill_2 FILLER_0_129_1075 ();
 sg13g2_fill_2 FILLER_0_129_1082 ();
 sg13g2_fill_4 FILLER_0_129_1092 ();
 sg13g2_fill_8 FILLER_0_129_1101 ();
 sg13g2_fill_8 FILLER_0_129_1109 ();
 sg13g2_fill_8 FILLER_0_129_1117 ();
 sg13g2_fill_8 FILLER_0_129_1125 ();
 sg13g2_fill_8 FILLER_0_129_1133 ();
 sg13g2_fill_2 FILLER_0_129_1141 ();
 sg13g2_fill_2 FILLER_0_129_1149 ();
 sg13g2_fill_1 FILLER_0_129_1151 ();
 sg13g2_fill_2 FILLER_0_129_1156 ();
 sg13g2_fill_1 FILLER_0_129_1158 ();
 sg13g2_fill_2 FILLER_0_129_1164 ();
 sg13g2_fill_1 FILLER_0_129_1166 ();
 sg13g2_fill_4 FILLER_0_129_1172 ();
 sg13g2_fill_1 FILLER_0_129_1176 ();
 sg13g2_fill_8 FILLER_0_129_1181 ();
 sg13g2_fill_8 FILLER_0_129_1189 ();
 sg13g2_fill_8 FILLER_0_129_1197 ();
 sg13g2_fill_4 FILLER_0_129_1205 ();
 sg13g2_fill_2 FILLER_0_129_1209 ();
 sg13g2_fill_1 FILLER_0_129_1211 ();
 sg13g2_fill_2 FILLER_0_129_1216 ();
 sg13g2_fill_2 FILLER_0_129_1223 ();
 sg13g2_fill_2 FILLER_0_129_1229 ();
 sg13g2_fill_2 FILLER_0_129_1236 ();
 sg13g2_fill_4 FILLER_0_129_1243 ();
 sg13g2_fill_1 FILLER_0_129_1247 ();
 sg13g2_fill_8 FILLER_0_129_1253 ();
 sg13g2_fill_1 FILLER_0_129_1261 ();
 sg13g2_fill_4 FILLER_0_129_1270 ();
 sg13g2_fill_2 FILLER_0_129_1274 ();
 sg13g2_fill_2 FILLER_0_129_1280 ();
 sg13g2_fill_8 FILLER_0_129_1288 ();
 sg13g2_fill_1 FILLER_0_129_1296 ();
 sg13g2_fill_8 FILLER_0_130_0 ();
 sg13g2_fill_8 FILLER_0_130_8 ();
 sg13g2_fill_8 FILLER_0_130_16 ();
 sg13g2_fill_8 FILLER_0_130_24 ();
 sg13g2_fill_8 FILLER_0_130_32 ();
 sg13g2_fill_8 FILLER_0_130_40 ();
 sg13g2_fill_8 FILLER_0_130_48 ();
 sg13g2_fill_8 FILLER_0_130_56 ();
 sg13g2_fill_8 FILLER_0_130_64 ();
 sg13g2_fill_8 FILLER_0_130_72 ();
 sg13g2_fill_8 FILLER_0_130_80 ();
 sg13g2_fill_8 FILLER_0_130_88 ();
 sg13g2_fill_8 FILLER_0_130_96 ();
 sg13g2_fill_8 FILLER_0_130_104 ();
 sg13g2_fill_8 FILLER_0_130_112 ();
 sg13g2_fill_8 FILLER_0_130_120 ();
 sg13g2_fill_8 FILLER_0_130_128 ();
 sg13g2_fill_8 FILLER_0_130_136 ();
 sg13g2_fill_8 FILLER_0_130_144 ();
 sg13g2_fill_8 FILLER_0_130_152 ();
 sg13g2_fill_8 FILLER_0_130_160 ();
 sg13g2_fill_8 FILLER_0_130_168 ();
 sg13g2_fill_8 FILLER_0_130_176 ();
 sg13g2_fill_8 FILLER_0_130_184 ();
 sg13g2_fill_8 FILLER_0_130_192 ();
 sg13g2_fill_8 FILLER_0_130_200 ();
 sg13g2_fill_8 FILLER_0_130_208 ();
 sg13g2_fill_8 FILLER_0_130_216 ();
 sg13g2_fill_8 FILLER_0_130_224 ();
 sg13g2_fill_8 FILLER_0_130_232 ();
 sg13g2_fill_8 FILLER_0_130_240 ();
 sg13g2_fill_8 FILLER_0_130_248 ();
 sg13g2_fill_4 FILLER_0_130_261 ();
 sg13g2_fill_8 FILLER_0_130_269 ();
 sg13g2_fill_4 FILLER_0_130_277 ();
 sg13g2_fill_2 FILLER_0_130_281 ();
 sg13g2_fill_1 FILLER_0_130_283 ();
 sg13g2_fill_4 FILLER_0_130_310 ();
 sg13g2_fill_1 FILLER_0_130_314 ();
 sg13g2_fill_2 FILLER_0_130_320 ();
 sg13g2_fill_8 FILLER_0_130_326 ();
 sg13g2_fill_8 FILLER_0_130_334 ();
 sg13g2_fill_2 FILLER_0_130_342 ();
 sg13g2_fill_4 FILLER_0_130_349 ();
 sg13g2_fill_2 FILLER_0_130_357 ();
 sg13g2_fill_1 FILLER_0_130_359 ();
 sg13g2_fill_2 FILLER_0_130_364 ();
 sg13g2_fill_2 FILLER_0_130_372 ();
 sg13g2_fill_1 FILLER_0_130_374 ();
 sg13g2_fill_8 FILLER_0_130_380 ();
 sg13g2_fill_8 FILLER_0_130_388 ();
 sg13g2_fill_8 FILLER_0_130_396 ();
 sg13g2_fill_2 FILLER_0_130_404 ();
 sg13g2_fill_2 FILLER_0_130_432 ();
 sg13g2_fill_2 FILLER_0_130_439 ();
 sg13g2_fill_4 FILLER_0_130_447 ();
 sg13g2_fill_2 FILLER_0_130_451 ();
 sg13g2_fill_8 FILLER_0_130_457 ();
 sg13g2_fill_8 FILLER_0_130_465 ();
 sg13g2_fill_2 FILLER_0_130_473 ();
 sg13g2_fill_2 FILLER_0_130_480 ();
 sg13g2_fill_2 FILLER_0_130_508 ();
 sg13g2_fill_4 FILLER_0_130_514 ();
 sg13g2_fill_1 FILLER_0_130_518 ();
 sg13g2_fill_2 FILLER_0_130_524 ();
 sg13g2_fill_2 FILLER_0_130_552 ();
 sg13g2_fill_4 FILLER_0_130_564 ();
 sg13g2_fill_8 FILLER_0_130_573 ();
 sg13g2_fill_2 FILLER_0_130_581 ();
 sg13g2_fill_1 FILLER_0_130_583 ();
 sg13g2_fill_8 FILLER_0_130_589 ();
 sg13g2_fill_1 FILLER_0_130_597 ();
 sg13g2_fill_8 FILLER_0_130_603 ();
 sg13g2_fill_4 FILLER_0_130_617 ();
 sg13g2_fill_4 FILLER_0_130_626 ();
 sg13g2_fill_2 FILLER_0_130_630 ();
 sg13g2_fill_1 FILLER_0_130_632 ();
 sg13g2_fill_8 FILLER_0_130_638 ();
 sg13g2_fill_2 FILLER_0_130_651 ();
 sg13g2_fill_2 FILLER_0_130_679 ();
 sg13g2_fill_8 FILLER_0_130_685 ();
 sg13g2_fill_4 FILLER_0_130_693 ();
 sg13g2_fill_8 FILLER_0_130_707 ();
 sg13g2_fill_8 FILLER_0_130_715 ();
 sg13g2_fill_8 FILLER_0_130_723 ();
 sg13g2_fill_8 FILLER_0_130_731 ();
 sg13g2_fill_8 FILLER_0_130_739 ();
 sg13g2_fill_8 FILLER_0_130_747 ();
 sg13g2_fill_8 FILLER_0_130_755 ();
 sg13g2_fill_8 FILLER_0_130_763 ();
 sg13g2_fill_4 FILLER_0_130_771 ();
 sg13g2_fill_8 FILLER_0_130_780 ();
 sg13g2_fill_8 FILLER_0_130_788 ();
 sg13g2_fill_4 FILLER_0_130_796 ();
 sg13g2_fill_2 FILLER_0_130_805 ();
 sg13g2_fill_2 FILLER_0_130_811 ();
 sg13g2_fill_8 FILLER_0_130_817 ();
 sg13g2_fill_8 FILLER_0_130_825 ();
 sg13g2_fill_8 FILLER_0_130_833 ();
 sg13g2_fill_8 FILLER_0_130_841 ();
 sg13g2_fill_4 FILLER_0_130_849 ();
 sg13g2_fill_1 FILLER_0_130_853 ();
 sg13g2_fill_4 FILLER_0_130_860 ();
 sg13g2_fill_2 FILLER_0_130_864 ();
 sg13g2_fill_1 FILLER_0_130_866 ();
 sg13g2_fill_4 FILLER_0_130_872 ();
 sg13g2_fill_1 FILLER_0_130_876 ();
 sg13g2_fill_2 FILLER_0_130_882 ();
 sg13g2_fill_2 FILLER_0_130_889 ();
 sg13g2_fill_2 FILLER_0_130_896 ();
 sg13g2_fill_8 FILLER_0_130_902 ();
 sg13g2_fill_4 FILLER_0_130_910 ();
 sg13g2_fill_2 FILLER_0_130_914 ();
 sg13g2_fill_1 FILLER_0_130_916 ();
 sg13g2_fill_4 FILLER_0_130_922 ();
 sg13g2_fill_1 FILLER_0_130_926 ();
 sg13g2_fill_2 FILLER_0_130_931 ();
 sg13g2_fill_1 FILLER_0_130_933 ();
 sg13g2_fill_4 FILLER_0_130_939 ();
 sg13g2_fill_4 FILLER_0_130_964 ();
 sg13g2_fill_4 FILLER_0_130_994 ();
 sg13g2_fill_8 FILLER_0_130_1003 ();
 sg13g2_fill_8 FILLER_0_130_1011 ();
 sg13g2_fill_8 FILLER_0_130_1019 ();
 sg13g2_fill_8 FILLER_0_130_1027 ();
 sg13g2_fill_8 FILLER_0_130_1035 ();
 sg13g2_fill_8 FILLER_0_130_1043 ();
 sg13g2_fill_8 FILLER_0_130_1051 ();
 sg13g2_fill_2 FILLER_0_130_1063 ();
 sg13g2_fill_8 FILLER_0_130_1070 ();
 sg13g2_fill_2 FILLER_0_130_1078 ();
 sg13g2_fill_1 FILLER_0_130_1080 ();
 sg13g2_fill_2 FILLER_0_130_1086 ();
 sg13g2_fill_2 FILLER_0_130_1096 ();
 sg13g2_fill_4 FILLER_0_130_1103 ();
 sg13g2_fill_1 FILLER_0_130_1107 ();
 sg13g2_fill_4 FILLER_0_130_1111 ();
 sg13g2_fill_1 FILLER_0_130_1115 ();
 sg13g2_fill_2 FILLER_0_130_1142 ();
 sg13g2_fill_2 FILLER_0_130_1149 ();
 sg13g2_fill_2 FILLER_0_130_1156 ();
 sg13g2_fill_1 FILLER_0_130_1158 ();
 sg13g2_fill_2 FILLER_0_130_1165 ();
 sg13g2_fill_1 FILLER_0_130_1167 ();
 sg13g2_fill_4 FILLER_0_130_1174 ();
 sg13g2_fill_4 FILLER_0_130_1186 ();
 sg13g2_fill_2 FILLER_0_130_1190 ();
 sg13g2_fill_4 FILLER_0_130_1197 ();
 sg13g2_fill_2 FILLER_0_130_1201 ();
 sg13g2_fill_1 FILLER_0_130_1203 ();
 sg13g2_fill_2 FILLER_0_130_1209 ();
 sg13g2_fill_8 FILLER_0_130_1219 ();
 sg13g2_fill_4 FILLER_0_130_1227 ();
 sg13g2_fill_1 FILLER_0_130_1231 ();
 sg13g2_fill_4 FILLER_0_130_1242 ();
 sg13g2_fill_2 FILLER_0_130_1246 ();
 sg13g2_fill_1 FILLER_0_130_1248 ();
 sg13g2_fill_2 FILLER_0_130_1275 ();
 sg13g2_fill_8 FILLER_0_130_1285 ();
 sg13g2_fill_4 FILLER_0_130_1293 ();
 sg13g2_fill_8 FILLER_0_131_0 ();
 sg13g2_fill_8 FILLER_0_131_8 ();
 sg13g2_fill_8 FILLER_0_131_16 ();
 sg13g2_fill_8 FILLER_0_131_24 ();
 sg13g2_fill_8 FILLER_0_131_32 ();
 sg13g2_fill_8 FILLER_0_131_40 ();
 sg13g2_fill_8 FILLER_0_131_48 ();
 sg13g2_fill_8 FILLER_0_131_56 ();
 sg13g2_fill_8 FILLER_0_131_64 ();
 sg13g2_fill_8 FILLER_0_131_72 ();
 sg13g2_fill_8 FILLER_0_131_80 ();
 sg13g2_fill_8 FILLER_0_131_88 ();
 sg13g2_fill_8 FILLER_0_131_96 ();
 sg13g2_fill_8 FILLER_0_131_104 ();
 sg13g2_fill_8 FILLER_0_131_112 ();
 sg13g2_fill_8 FILLER_0_131_120 ();
 sg13g2_fill_8 FILLER_0_131_128 ();
 sg13g2_fill_8 FILLER_0_131_136 ();
 sg13g2_fill_8 FILLER_0_131_144 ();
 sg13g2_fill_8 FILLER_0_131_152 ();
 sg13g2_fill_8 FILLER_0_131_160 ();
 sg13g2_fill_8 FILLER_0_131_168 ();
 sg13g2_fill_8 FILLER_0_131_176 ();
 sg13g2_fill_8 FILLER_0_131_184 ();
 sg13g2_fill_8 FILLER_0_131_192 ();
 sg13g2_fill_8 FILLER_0_131_200 ();
 sg13g2_fill_8 FILLER_0_131_208 ();
 sg13g2_fill_8 FILLER_0_131_216 ();
 sg13g2_fill_8 FILLER_0_131_224 ();
 sg13g2_fill_8 FILLER_0_131_232 ();
 sg13g2_fill_8 FILLER_0_131_240 ();
 sg13g2_fill_4 FILLER_0_131_248 ();
 sg13g2_fill_4 FILLER_0_131_278 ();
 sg13g2_fill_2 FILLER_0_131_282 ();
 sg13g2_fill_2 FILLER_0_131_289 ();
 sg13g2_fill_2 FILLER_0_131_301 ();
 sg13g2_fill_2 FILLER_0_131_329 ();
 sg13g2_fill_8 FILLER_0_131_336 ();
 sg13g2_fill_1 FILLER_0_131_344 ();
 sg13g2_fill_4 FILLER_0_131_349 ();
 sg13g2_fill_2 FILLER_0_131_353 ();
 sg13g2_fill_1 FILLER_0_131_355 ();
 sg13g2_fill_8 FILLER_0_131_361 ();
 sg13g2_fill_8 FILLER_0_131_369 ();
 sg13g2_fill_8 FILLER_0_131_377 ();
 sg13g2_fill_8 FILLER_0_131_385 ();
 sg13g2_fill_8 FILLER_0_131_393 ();
 sg13g2_fill_4 FILLER_0_131_401 ();
 sg13g2_fill_2 FILLER_0_131_405 ();
 sg13g2_fill_1 FILLER_0_131_407 ();
 sg13g2_fill_2 FILLER_0_131_413 ();
 sg13g2_fill_4 FILLER_0_131_419 ();
 sg13g2_fill_2 FILLER_0_131_423 ();
 sg13g2_fill_2 FILLER_0_131_430 ();
 sg13g2_fill_2 FILLER_0_131_436 ();
 sg13g2_fill_2 FILLER_0_131_464 ();
 sg13g2_fill_1 FILLER_0_131_466 ();
 sg13g2_fill_4 FILLER_0_131_493 ();
 sg13g2_fill_2 FILLER_0_131_497 ();
 sg13g2_fill_1 FILLER_0_131_499 ();
 sg13g2_fill_8 FILLER_0_131_506 ();
 sg13g2_fill_8 FILLER_0_131_514 ();
 sg13g2_fill_8 FILLER_0_131_527 ();
 sg13g2_fill_2 FILLER_0_131_535 ();
 sg13g2_fill_8 FILLER_0_131_541 ();
 sg13g2_fill_8 FILLER_0_131_549 ();
 sg13g2_fill_1 FILLER_0_131_557 ();
 sg13g2_fill_8 FILLER_0_131_563 ();
 sg13g2_fill_2 FILLER_0_131_571 ();
 sg13g2_fill_2 FILLER_0_131_578 ();
 sg13g2_fill_8 FILLER_0_131_584 ();
 sg13g2_fill_8 FILLER_0_131_592 ();
 sg13g2_fill_4 FILLER_0_131_600 ();
 sg13g2_fill_2 FILLER_0_131_604 ();
 sg13g2_fill_2 FILLER_0_131_611 ();
 sg13g2_fill_8 FILLER_0_131_639 ();
 sg13g2_fill_8 FILLER_0_131_647 ();
 sg13g2_fill_8 FILLER_0_131_655 ();
 sg13g2_fill_8 FILLER_0_131_663 ();
 sg13g2_fill_2 FILLER_0_131_671 ();
 sg13g2_fill_1 FILLER_0_131_673 ();
 sg13g2_fill_2 FILLER_0_131_679 ();
 sg13g2_fill_2 FILLER_0_131_707 ();
 sg13g2_fill_8 FILLER_0_131_713 ();
 sg13g2_fill_2 FILLER_0_131_721 ();
 sg13g2_fill_8 FILLER_0_131_731 ();
 sg13g2_fill_8 FILLER_0_131_739 ();
 sg13g2_fill_8 FILLER_0_131_747 ();
 sg13g2_fill_8 FILLER_0_131_755 ();
 sg13g2_fill_8 FILLER_0_131_763 ();
 sg13g2_fill_8 FILLER_0_131_771 ();
 sg13g2_fill_4 FILLER_0_131_779 ();
 sg13g2_fill_2 FILLER_0_131_788 ();
 sg13g2_fill_1 FILLER_0_131_790 ();
 sg13g2_fill_4 FILLER_0_131_795 ();
 sg13g2_fill_2 FILLER_0_131_799 ();
 sg13g2_fill_1 FILLER_0_131_801 ();
 sg13g2_fill_8 FILLER_0_131_807 ();
 sg13g2_fill_8 FILLER_0_131_815 ();
 sg13g2_fill_8 FILLER_0_131_823 ();
 sg13g2_fill_1 FILLER_0_131_831 ();
 sg13g2_fill_4 FILLER_0_131_837 ();
 sg13g2_fill_1 FILLER_0_131_841 ();
 sg13g2_fill_2 FILLER_0_131_847 ();
 sg13g2_fill_1 FILLER_0_131_849 ();
 sg13g2_fill_4 FILLER_0_131_855 ();
 sg13g2_fill_2 FILLER_0_131_859 ();
 sg13g2_fill_4 FILLER_0_131_887 ();
 sg13g2_fill_2 FILLER_0_131_891 ();
 sg13g2_fill_8 FILLER_0_131_898 ();
 sg13g2_fill_8 FILLER_0_131_906 ();
 sg13g2_fill_2 FILLER_0_131_914 ();
 sg13g2_fill_2 FILLER_0_131_920 ();
 sg13g2_fill_2 FILLER_0_131_948 ();
 sg13g2_fill_2 FILLER_0_131_955 ();
 sg13g2_fill_2 FILLER_0_131_961 ();
 sg13g2_fill_2 FILLER_0_131_989 ();
 sg13g2_fill_2 FILLER_0_131_997 ();
 sg13g2_fill_1 FILLER_0_131_999 ();
 sg13g2_fill_4 FILLER_0_131_1005 ();
 sg13g2_fill_2 FILLER_0_131_1016 ();
 sg13g2_fill_4 FILLER_0_131_1023 ();
 sg13g2_fill_2 FILLER_0_131_1027 ();
 sg13g2_fill_8 FILLER_0_131_1035 ();
 sg13g2_fill_8 FILLER_0_131_1043 ();
 sg13g2_fill_2 FILLER_0_131_1051 ();
 sg13g2_fill_1 FILLER_0_131_1053 ();
 sg13g2_fill_2 FILLER_0_131_1058 ();
 sg13g2_fill_2 FILLER_0_131_1065 ();
 sg13g2_fill_8 FILLER_0_131_1072 ();
 sg13g2_fill_8 FILLER_0_131_1080 ();
 sg13g2_fill_1 FILLER_0_131_1088 ();
 sg13g2_fill_2 FILLER_0_131_1097 ();
 sg13g2_fill_2 FILLER_0_131_1103 ();
 sg13g2_fill_4 FILLER_0_131_1109 ();
 sg13g2_fill_1 FILLER_0_131_1113 ();
 sg13g2_fill_2 FILLER_0_131_1124 ();
 sg13g2_fill_4 FILLER_0_131_1136 ();
 sg13g2_fill_4 FILLER_0_131_1148 ();
 sg13g2_fill_1 FILLER_0_131_1152 ();
 sg13g2_fill_2 FILLER_0_131_1159 ();
 sg13g2_fill_2 FILLER_0_131_1166 ();
 sg13g2_fill_1 FILLER_0_131_1168 ();
 sg13g2_fill_8 FILLER_0_131_1174 ();
 sg13g2_fill_4 FILLER_0_131_1182 ();
 sg13g2_fill_2 FILLER_0_131_1194 ();
 sg13g2_fill_1 FILLER_0_131_1196 ();
 sg13g2_fill_2 FILLER_0_131_1202 ();
 sg13g2_fill_4 FILLER_0_131_1208 ();
 sg13g2_fill_2 FILLER_0_131_1218 ();
 sg13g2_fill_2 FILLER_0_131_1225 ();
 sg13g2_fill_8 FILLER_0_131_1232 ();
 sg13g2_fill_8 FILLER_0_131_1240 ();
 sg13g2_fill_4 FILLER_0_131_1248 ();
 sg13g2_fill_1 FILLER_0_131_1252 ();
 sg13g2_fill_2 FILLER_0_131_1263 ();
 sg13g2_fill_8 FILLER_0_131_1275 ();
 sg13g2_fill_8 FILLER_0_131_1287 ();
 sg13g2_fill_2 FILLER_0_131_1295 ();
 sg13g2_fill_8 FILLER_0_132_0 ();
 sg13g2_fill_8 FILLER_0_132_8 ();
 sg13g2_fill_8 FILLER_0_132_16 ();
 sg13g2_fill_8 FILLER_0_132_24 ();
 sg13g2_fill_8 FILLER_0_132_32 ();
 sg13g2_fill_8 FILLER_0_132_40 ();
 sg13g2_fill_8 FILLER_0_132_48 ();
 sg13g2_fill_8 FILLER_0_132_56 ();
 sg13g2_fill_8 FILLER_0_132_64 ();
 sg13g2_fill_8 FILLER_0_132_72 ();
 sg13g2_fill_8 FILLER_0_132_80 ();
 sg13g2_fill_8 FILLER_0_132_88 ();
 sg13g2_fill_8 FILLER_0_132_96 ();
 sg13g2_fill_8 FILLER_0_132_104 ();
 sg13g2_fill_8 FILLER_0_132_112 ();
 sg13g2_fill_8 FILLER_0_132_120 ();
 sg13g2_fill_8 FILLER_0_132_128 ();
 sg13g2_fill_8 FILLER_0_132_136 ();
 sg13g2_fill_8 FILLER_0_132_144 ();
 sg13g2_fill_8 FILLER_0_132_152 ();
 sg13g2_fill_8 FILLER_0_132_160 ();
 sg13g2_fill_8 FILLER_0_132_168 ();
 sg13g2_fill_8 FILLER_0_132_176 ();
 sg13g2_fill_8 FILLER_0_132_184 ();
 sg13g2_fill_8 FILLER_0_132_192 ();
 sg13g2_fill_8 FILLER_0_132_200 ();
 sg13g2_fill_8 FILLER_0_132_208 ();
 sg13g2_fill_8 FILLER_0_132_216 ();
 sg13g2_fill_8 FILLER_0_132_224 ();
 sg13g2_fill_8 FILLER_0_132_232 ();
 sg13g2_fill_8 FILLER_0_132_240 ();
 sg13g2_fill_8 FILLER_0_132_248 ();
 sg13g2_fill_8 FILLER_0_132_256 ();
 sg13g2_fill_1 FILLER_0_132_264 ();
 sg13g2_fill_4 FILLER_0_132_291 ();
 sg13g2_fill_1 FILLER_0_132_295 ();
 sg13g2_fill_8 FILLER_0_132_317 ();
 sg13g2_fill_8 FILLER_0_132_325 ();
 sg13g2_fill_8 FILLER_0_132_333 ();
 sg13g2_fill_8 FILLER_0_132_341 ();
 sg13g2_fill_8 FILLER_0_132_349 ();
 sg13g2_fill_8 FILLER_0_132_357 ();
 sg13g2_fill_8 FILLER_0_132_365 ();
 sg13g2_fill_8 FILLER_0_132_373 ();
 sg13g2_fill_2 FILLER_0_132_381 ();
 sg13g2_fill_1 FILLER_0_132_383 ();
 sg13g2_fill_2 FILLER_0_132_389 ();
 sg13g2_fill_8 FILLER_0_132_417 ();
 sg13g2_fill_4 FILLER_0_132_425 ();
 sg13g2_fill_2 FILLER_0_132_429 ();
 sg13g2_fill_1 FILLER_0_132_431 ();
 sg13g2_fill_8 FILLER_0_132_437 ();
 sg13g2_fill_8 FILLER_0_132_445 ();
 sg13g2_fill_8 FILLER_0_132_453 ();
 sg13g2_fill_8 FILLER_0_132_461 ();
 sg13g2_fill_8 FILLER_0_132_469 ();
 sg13g2_fill_2 FILLER_0_132_482 ();
 sg13g2_fill_4 FILLER_0_132_488 ();
 sg13g2_fill_2 FILLER_0_132_492 ();
 sg13g2_fill_1 FILLER_0_132_494 ();
 sg13g2_fill_8 FILLER_0_132_500 ();
 sg13g2_fill_8 FILLER_0_132_508 ();
 sg13g2_fill_8 FILLER_0_132_516 ();
 sg13g2_fill_8 FILLER_0_132_524 ();
 sg13g2_fill_8 FILLER_0_132_532 ();
 sg13g2_fill_8 FILLER_0_132_540 ();
 sg13g2_fill_4 FILLER_0_132_548 ();
 sg13g2_fill_8 FILLER_0_132_557 ();
 sg13g2_fill_4 FILLER_0_132_565 ();
 sg13g2_fill_2 FILLER_0_132_569 ();
 sg13g2_fill_2 FILLER_0_132_597 ();
 sg13g2_fill_4 FILLER_0_132_603 ();
 sg13g2_fill_2 FILLER_0_132_607 ();
 sg13g2_fill_1 FILLER_0_132_609 ();
 sg13g2_fill_2 FILLER_0_132_615 ();
 sg13g2_fill_2 FILLER_0_132_622 ();
 sg13g2_fill_4 FILLER_0_132_628 ();
 sg13g2_fill_1 FILLER_0_132_632 ();
 sg13g2_fill_2 FILLER_0_132_637 ();
 sg13g2_fill_1 FILLER_0_132_639 ();
 sg13g2_fill_8 FILLER_0_132_645 ();
 sg13g2_fill_8 FILLER_0_132_653 ();
 sg13g2_fill_8 FILLER_0_132_661 ();
 sg13g2_fill_8 FILLER_0_132_669 ();
 sg13g2_fill_8 FILLER_0_132_677 ();
 sg13g2_fill_8 FILLER_0_132_685 ();
 sg13g2_fill_4 FILLER_0_132_693 ();
 sg13g2_fill_8 FILLER_0_132_705 ();
 sg13g2_fill_8 FILLER_0_132_713 ();
 sg13g2_fill_8 FILLER_0_132_721 ();
 sg13g2_fill_8 FILLER_0_132_729 ();
 sg13g2_fill_2 FILLER_0_132_743 ();
 sg13g2_fill_2 FILLER_0_132_751 ();
 sg13g2_fill_1 FILLER_0_132_753 ();
 sg13g2_fill_8 FILLER_0_132_759 ();
 sg13g2_fill_2 FILLER_0_132_767 ();
 sg13g2_fill_2 FILLER_0_132_773 ();
 sg13g2_fill_8 FILLER_0_132_801 ();
 sg13g2_fill_8 FILLER_0_132_809 ();
 sg13g2_fill_2 FILLER_0_132_817 ();
 sg13g2_fill_4 FILLER_0_132_824 ();
 sg13g2_fill_1 FILLER_0_132_828 ();
 sg13g2_fill_8 FILLER_0_132_833 ();
 sg13g2_fill_4 FILLER_0_132_841 ();
 sg13g2_fill_2 FILLER_0_132_845 ();
 sg13g2_fill_1 FILLER_0_132_847 ();
 sg13g2_fill_4 FILLER_0_132_853 ();
 sg13g2_fill_2 FILLER_0_132_862 ();
 sg13g2_fill_8 FILLER_0_132_868 ();
 sg13g2_fill_8 FILLER_0_132_876 ();
 sg13g2_fill_8 FILLER_0_132_884 ();
 sg13g2_fill_2 FILLER_0_132_892 ();
 sg13g2_fill_4 FILLER_0_132_900 ();
 sg13g2_fill_2 FILLER_0_132_904 ();
 sg13g2_fill_1 FILLER_0_132_906 ();
 sg13g2_fill_8 FILLER_0_132_916 ();
 sg13g2_fill_8 FILLER_0_132_924 ();
 sg13g2_fill_8 FILLER_0_132_932 ();
 sg13g2_fill_2 FILLER_0_132_940 ();
 sg13g2_fill_1 FILLER_0_132_942 ();
 sg13g2_fill_2 FILLER_0_132_947 ();
 sg13g2_fill_1 FILLER_0_132_949 ();
 sg13g2_fill_4 FILLER_0_132_955 ();
 sg13g2_fill_2 FILLER_0_132_959 ();
 sg13g2_fill_2 FILLER_0_132_966 ();
 sg13g2_fill_1 FILLER_0_132_968 ();
 sg13g2_fill_8 FILLER_0_132_976 ();
 sg13g2_fill_8 FILLER_0_132_984 ();
 sg13g2_fill_4 FILLER_0_132_992 ();
 sg13g2_fill_2 FILLER_0_132_996 ();
 sg13g2_fill_1 FILLER_0_132_998 ();
 sg13g2_fill_8 FILLER_0_132_1003 ();
 sg13g2_fill_8 FILLER_0_132_1011 ();
 sg13g2_fill_8 FILLER_0_132_1019 ();
 sg13g2_fill_2 FILLER_0_132_1027 ();
 sg13g2_fill_1 FILLER_0_132_1029 ();
 sg13g2_fill_2 FILLER_0_132_1037 ();
 sg13g2_fill_8 FILLER_0_132_1044 ();
 sg13g2_fill_8 FILLER_0_132_1052 ();
 sg13g2_fill_8 FILLER_0_132_1060 ();
 sg13g2_fill_8 FILLER_0_132_1068 ();
 sg13g2_fill_8 FILLER_0_132_1076 ();
 sg13g2_fill_8 FILLER_0_132_1084 ();
 sg13g2_fill_8 FILLER_0_132_1092 ();
 sg13g2_fill_8 FILLER_0_132_1100 ();
 sg13g2_fill_8 FILLER_0_132_1108 ();
 sg13g2_fill_8 FILLER_0_132_1116 ();
 sg13g2_fill_8 FILLER_0_132_1124 ();
 sg13g2_fill_8 FILLER_0_132_1132 ();
 sg13g2_fill_8 FILLER_0_132_1140 ();
 sg13g2_fill_8 FILLER_0_132_1148 ();
 sg13g2_fill_8 FILLER_0_132_1156 ();
 sg13g2_fill_2 FILLER_0_132_1164 ();
 sg13g2_fill_1 FILLER_0_132_1166 ();
 sg13g2_fill_2 FILLER_0_132_1171 ();
 sg13g2_fill_8 FILLER_0_132_1177 ();
 sg13g2_fill_2 FILLER_0_132_1193 ();
 sg13g2_fill_2 FILLER_0_132_1200 ();
 sg13g2_fill_2 FILLER_0_132_1210 ();
 sg13g2_fill_2 FILLER_0_132_1216 ();
 sg13g2_fill_1 FILLER_0_132_1218 ();
 sg13g2_fill_4 FILLER_0_132_1224 ();
 sg13g2_fill_2 FILLER_0_132_1233 ();
 sg13g2_fill_8 FILLER_0_132_1238 ();
 sg13g2_fill_1 FILLER_0_132_1246 ();
 sg13g2_fill_8 FILLER_0_132_1252 ();
 sg13g2_fill_4 FILLER_0_132_1260 ();
 sg13g2_fill_1 FILLER_0_132_1264 ();
 sg13g2_fill_8 FILLER_0_132_1269 ();
 sg13g2_fill_8 FILLER_0_132_1277 ();
 sg13g2_fill_8 FILLER_0_132_1285 ();
 sg13g2_fill_4 FILLER_0_132_1293 ();
 sg13g2_fill_8 FILLER_0_133_0 ();
 sg13g2_fill_8 FILLER_0_133_8 ();
 sg13g2_fill_8 FILLER_0_133_16 ();
 sg13g2_fill_8 FILLER_0_133_24 ();
 sg13g2_fill_8 FILLER_0_133_32 ();
 sg13g2_fill_8 FILLER_0_133_40 ();
 sg13g2_fill_8 FILLER_0_133_48 ();
 sg13g2_fill_8 FILLER_0_133_56 ();
 sg13g2_fill_8 FILLER_0_133_64 ();
 sg13g2_fill_8 FILLER_0_133_72 ();
 sg13g2_fill_8 FILLER_0_133_80 ();
 sg13g2_fill_8 FILLER_0_133_88 ();
 sg13g2_fill_8 FILLER_0_133_96 ();
 sg13g2_fill_8 FILLER_0_133_104 ();
 sg13g2_fill_8 FILLER_0_133_112 ();
 sg13g2_fill_8 FILLER_0_133_120 ();
 sg13g2_fill_8 FILLER_0_133_128 ();
 sg13g2_fill_8 FILLER_0_133_136 ();
 sg13g2_fill_8 FILLER_0_133_144 ();
 sg13g2_fill_8 FILLER_0_133_152 ();
 sg13g2_fill_8 FILLER_0_133_160 ();
 sg13g2_fill_8 FILLER_0_133_168 ();
 sg13g2_fill_8 FILLER_0_133_176 ();
 sg13g2_fill_8 FILLER_0_133_184 ();
 sg13g2_fill_8 FILLER_0_133_192 ();
 sg13g2_fill_8 FILLER_0_133_200 ();
 sg13g2_fill_8 FILLER_0_133_208 ();
 sg13g2_fill_8 FILLER_0_133_216 ();
 sg13g2_fill_8 FILLER_0_133_224 ();
 sg13g2_fill_8 FILLER_0_133_232 ();
 sg13g2_fill_8 FILLER_0_133_240 ();
 sg13g2_fill_8 FILLER_0_133_248 ();
 sg13g2_fill_8 FILLER_0_133_256 ();
 sg13g2_fill_8 FILLER_0_133_264 ();
 sg13g2_fill_8 FILLER_0_133_272 ();
 sg13g2_fill_1 FILLER_0_133_280 ();
 sg13g2_fill_8 FILLER_0_133_285 ();
 sg13g2_fill_8 FILLER_0_133_293 ();
 sg13g2_fill_8 FILLER_0_133_301 ();
 sg13g2_fill_8 FILLER_0_133_309 ();
 sg13g2_fill_2 FILLER_0_133_317 ();
 sg13g2_fill_1 FILLER_0_133_319 ();
 sg13g2_fill_8 FILLER_0_133_324 ();
 sg13g2_fill_8 FILLER_0_133_332 ();
 sg13g2_fill_4 FILLER_0_133_340 ();
 sg13g2_fill_1 FILLER_0_133_344 ();
 sg13g2_fill_2 FILLER_0_133_350 ();
 sg13g2_fill_8 FILLER_0_133_356 ();
 sg13g2_fill_8 FILLER_0_133_364 ();
 sg13g2_fill_2 FILLER_0_133_372 ();
 sg13g2_fill_8 FILLER_0_133_381 ();
 sg13g2_fill_8 FILLER_0_133_389 ();
 sg13g2_fill_8 FILLER_0_133_397 ();
 sg13g2_fill_8 FILLER_0_133_405 ();
 sg13g2_fill_4 FILLER_0_133_413 ();
 sg13g2_fill_2 FILLER_0_133_417 ();
 sg13g2_fill_4 FILLER_0_133_423 ();
 sg13g2_fill_2 FILLER_0_133_427 ();
 sg13g2_fill_8 FILLER_0_133_435 ();
 sg13g2_fill_8 FILLER_0_133_443 ();
 sg13g2_fill_8 FILLER_0_133_451 ();
 sg13g2_fill_8 FILLER_0_133_459 ();
 sg13g2_fill_8 FILLER_0_133_467 ();
 sg13g2_fill_8 FILLER_0_133_475 ();
 sg13g2_fill_8 FILLER_0_133_483 ();
 sg13g2_fill_4 FILLER_0_133_491 ();
 sg13g2_fill_1 FILLER_0_133_495 ();
 sg13g2_fill_4 FILLER_0_133_501 ();
 sg13g2_fill_4 FILLER_0_133_510 ();
 sg13g2_fill_1 FILLER_0_133_514 ();
 sg13g2_fill_8 FILLER_0_133_519 ();
 sg13g2_fill_8 FILLER_0_133_527 ();
 sg13g2_fill_8 FILLER_0_133_535 ();
 sg13g2_fill_8 FILLER_0_133_543 ();
 sg13g2_fill_8 FILLER_0_133_551 ();
 sg13g2_fill_8 FILLER_0_133_559 ();
 sg13g2_fill_4 FILLER_0_133_567 ();
 sg13g2_fill_1 FILLER_0_133_571 ();
 sg13g2_fill_8 FILLER_0_133_577 ();
 sg13g2_fill_8 FILLER_0_133_585 ();
 sg13g2_fill_8 FILLER_0_133_593 ();
 sg13g2_fill_8 FILLER_0_133_601 ();
 sg13g2_fill_8 FILLER_0_133_609 ();
 sg13g2_fill_8 FILLER_0_133_617 ();
 sg13g2_fill_8 FILLER_0_133_625 ();
 sg13g2_fill_8 FILLER_0_133_633 ();
 sg13g2_fill_2 FILLER_0_133_641 ();
 sg13g2_fill_1 FILLER_0_133_643 ();
 sg13g2_fill_4 FILLER_0_133_649 ();
 sg13g2_fill_2 FILLER_0_133_657 ();
 sg13g2_fill_2 FILLER_0_133_664 ();
 sg13g2_fill_2 FILLER_0_133_671 ();
 sg13g2_fill_8 FILLER_0_133_678 ();
 sg13g2_fill_2 FILLER_0_133_686 ();
 sg13g2_fill_1 FILLER_0_133_688 ();
 sg13g2_fill_8 FILLER_0_133_694 ();
 sg13g2_fill_8 FILLER_0_133_702 ();
 sg13g2_fill_8 FILLER_0_133_710 ();
 sg13g2_fill_1 FILLER_0_133_718 ();
 sg13g2_fill_2 FILLER_0_133_724 ();
 sg13g2_fill_2 FILLER_0_133_730 ();
 sg13g2_fill_4 FILLER_0_133_737 ();
 sg13g2_fill_2 FILLER_0_133_741 ();
 sg13g2_fill_2 FILLER_0_133_769 ();
 sg13g2_fill_8 FILLER_0_133_792 ();
 sg13g2_fill_4 FILLER_0_133_800 ();
 sg13g2_fill_2 FILLER_0_133_804 ();
 sg13g2_fill_1 FILLER_0_133_806 ();
 sg13g2_fill_2 FILLER_0_133_812 ();
 sg13g2_fill_2 FILLER_0_133_818 ();
 sg13g2_fill_2 FILLER_0_133_846 ();
 sg13g2_fill_8 FILLER_0_133_853 ();
 sg13g2_fill_8 FILLER_0_133_861 ();
 sg13g2_fill_8 FILLER_0_133_869 ();
 sg13g2_fill_1 FILLER_0_133_877 ();
 sg13g2_fill_8 FILLER_0_133_904 ();
 sg13g2_fill_4 FILLER_0_133_912 ();
 sg13g2_fill_2 FILLER_0_133_924 ();
 sg13g2_fill_1 FILLER_0_133_926 ();
 sg13g2_fill_2 FILLER_0_133_932 ();
 sg13g2_fill_8 FILLER_0_133_938 ();
 sg13g2_fill_8 FILLER_0_133_946 ();
 sg13g2_fill_8 FILLER_0_133_954 ();
 sg13g2_fill_4 FILLER_0_133_962 ();
 sg13g2_fill_8 FILLER_0_133_978 ();
 sg13g2_fill_8 FILLER_0_133_986 ();
 sg13g2_fill_4 FILLER_0_133_994 ();
 sg13g2_fill_1 FILLER_0_133_998 ();
 sg13g2_fill_8 FILLER_0_133_1007 ();
 sg13g2_fill_8 FILLER_0_133_1015 ();
 sg13g2_fill_8 FILLER_0_133_1023 ();
 sg13g2_fill_4 FILLER_0_133_1031 ();
 sg13g2_fill_4 FILLER_0_133_1043 ();
 sg13g2_fill_2 FILLER_0_133_1047 ();
 sg13g2_fill_1 FILLER_0_133_1049 ();
 sg13g2_fill_8 FILLER_0_133_1055 ();
 sg13g2_fill_4 FILLER_0_133_1063 ();
 sg13g2_fill_1 FILLER_0_133_1067 ();
 sg13g2_fill_8 FILLER_0_133_1073 ();
 sg13g2_fill_2 FILLER_0_133_1081 ();
 sg13g2_fill_1 FILLER_0_133_1083 ();
 sg13g2_fill_8 FILLER_0_133_1088 ();
 sg13g2_fill_8 FILLER_0_133_1096 ();
 sg13g2_fill_8 FILLER_0_133_1104 ();
 sg13g2_fill_8 FILLER_0_133_1112 ();
 sg13g2_fill_4 FILLER_0_133_1120 ();
 sg13g2_fill_8 FILLER_0_133_1129 ();
 sg13g2_fill_2 FILLER_0_133_1137 ();
 sg13g2_fill_1 FILLER_0_133_1139 ();
 sg13g2_fill_8 FILLER_0_133_1144 ();
 sg13g2_fill_8 FILLER_0_133_1152 ();
 sg13g2_fill_8 FILLER_0_133_1160 ();
 sg13g2_fill_8 FILLER_0_133_1168 ();
 sg13g2_fill_8 FILLER_0_133_1176 ();
 sg13g2_fill_4 FILLER_0_133_1184 ();
 sg13g2_fill_1 FILLER_0_133_1188 ();
 sg13g2_fill_4 FILLER_0_133_1196 ();
 sg13g2_fill_8 FILLER_0_133_1207 ();
 sg13g2_fill_8 FILLER_0_133_1215 ();
 sg13g2_fill_4 FILLER_0_133_1223 ();
 sg13g2_fill_2 FILLER_0_133_1227 ();
 sg13g2_fill_8 FILLER_0_133_1233 ();
 sg13g2_fill_8 FILLER_0_133_1241 ();
 sg13g2_fill_8 FILLER_0_133_1249 ();
 sg13g2_fill_8 FILLER_0_133_1257 ();
 sg13g2_fill_2 FILLER_0_133_1265 ();
 sg13g2_fill_8 FILLER_0_133_1270 ();
 sg13g2_fill_8 FILLER_0_133_1278 ();
 sg13g2_fill_8 FILLER_0_133_1286 ();
 sg13g2_fill_2 FILLER_0_133_1294 ();
 sg13g2_fill_1 FILLER_0_133_1296 ();
 sg13g2_fill_8 FILLER_0_134_0 ();
 sg13g2_fill_8 FILLER_0_134_8 ();
 sg13g2_fill_8 FILLER_0_134_16 ();
 sg13g2_fill_8 FILLER_0_134_24 ();
 sg13g2_fill_8 FILLER_0_134_32 ();
 sg13g2_fill_8 FILLER_0_134_40 ();
 sg13g2_fill_8 FILLER_0_134_48 ();
 sg13g2_fill_8 FILLER_0_134_56 ();
 sg13g2_fill_8 FILLER_0_134_64 ();
 sg13g2_fill_8 FILLER_0_134_72 ();
 sg13g2_fill_8 FILLER_0_134_80 ();
 sg13g2_fill_8 FILLER_0_134_88 ();
 sg13g2_fill_8 FILLER_0_134_96 ();
 sg13g2_fill_8 FILLER_0_134_104 ();
 sg13g2_fill_8 FILLER_0_134_112 ();
 sg13g2_fill_8 FILLER_0_134_120 ();
 sg13g2_fill_8 FILLER_0_134_128 ();
 sg13g2_fill_8 FILLER_0_134_136 ();
 sg13g2_fill_8 FILLER_0_134_144 ();
 sg13g2_fill_8 FILLER_0_134_152 ();
 sg13g2_fill_8 FILLER_0_134_160 ();
 sg13g2_fill_8 FILLER_0_134_168 ();
 sg13g2_fill_8 FILLER_0_134_176 ();
 sg13g2_fill_8 FILLER_0_134_184 ();
 sg13g2_fill_8 FILLER_0_134_192 ();
 sg13g2_fill_8 FILLER_0_134_200 ();
 sg13g2_fill_8 FILLER_0_134_208 ();
 sg13g2_fill_8 FILLER_0_134_216 ();
 sg13g2_fill_8 FILLER_0_134_224 ();
 sg13g2_fill_8 FILLER_0_134_232 ();
 sg13g2_fill_8 FILLER_0_134_240 ();
 sg13g2_fill_8 FILLER_0_134_248 ();
 sg13g2_fill_8 FILLER_0_134_256 ();
 sg13g2_fill_2 FILLER_0_134_264 ();
 sg13g2_fill_1 FILLER_0_134_266 ();
 sg13g2_fill_8 FILLER_0_134_272 ();
 sg13g2_fill_8 FILLER_0_134_280 ();
 sg13g2_fill_8 FILLER_0_134_288 ();
 sg13g2_fill_4 FILLER_0_134_296 ();
 sg13g2_fill_2 FILLER_0_134_300 ();
 sg13g2_fill_8 FILLER_0_134_307 ();
 sg13g2_fill_8 FILLER_0_134_319 ();
 sg13g2_fill_8 FILLER_0_134_327 ();
 sg13g2_fill_4 FILLER_0_134_335 ();
 sg13g2_fill_1 FILLER_0_134_339 ();
 sg13g2_fill_8 FILLER_0_134_366 ();
 sg13g2_fill_8 FILLER_0_134_374 ();
 sg13g2_fill_8 FILLER_0_134_382 ();
 sg13g2_fill_4 FILLER_0_134_390 ();
 sg13g2_fill_2 FILLER_0_134_400 ();
 sg13g2_fill_4 FILLER_0_134_428 ();
 sg13g2_fill_2 FILLER_0_134_439 ();
 sg13g2_fill_8 FILLER_0_134_446 ();
 sg13g2_fill_8 FILLER_0_134_454 ();
 sg13g2_fill_1 FILLER_0_134_462 ();
 sg13g2_fill_4 FILLER_0_134_468 ();
 sg13g2_fill_2 FILLER_0_134_476 ();
 sg13g2_fill_4 FILLER_0_134_483 ();
 sg13g2_fill_8 FILLER_0_134_491 ();
 sg13g2_fill_2 FILLER_0_134_499 ();
 sg13g2_fill_4 FILLER_0_134_527 ();
 sg13g2_fill_2 FILLER_0_134_531 ();
 sg13g2_fill_2 FILLER_0_134_554 ();
 sg13g2_fill_1 FILLER_0_134_556 ();
 sg13g2_fill_4 FILLER_0_134_567 ();
 sg13g2_fill_2 FILLER_0_134_571 ();
 sg13g2_fill_4 FILLER_0_134_581 ();
 sg13g2_fill_1 FILLER_0_134_585 ();
 sg13g2_fill_2 FILLER_0_134_592 ();
 sg13g2_fill_2 FILLER_0_134_602 ();
 sg13g2_fill_2 FILLER_0_134_609 ();
 sg13g2_fill_4 FILLER_0_134_618 ();
 sg13g2_fill_2 FILLER_0_134_627 ();
 sg13g2_fill_1 FILLER_0_134_629 ();
 sg13g2_fill_4 FILLER_0_134_634 ();
 sg13g2_fill_2 FILLER_0_134_638 ();
 sg13g2_fill_1 FILLER_0_134_640 ();
 sg13g2_fill_2 FILLER_0_134_667 ();
 sg13g2_fill_4 FILLER_0_134_675 ();
 sg13g2_fill_2 FILLER_0_134_679 ();
 sg13g2_fill_2 FILLER_0_134_689 ();
 sg13g2_fill_2 FILLER_0_134_696 ();
 sg13g2_fill_8 FILLER_0_134_724 ();
 sg13g2_fill_8 FILLER_0_134_732 ();
 sg13g2_fill_4 FILLER_0_134_740 ();
 sg13g2_fill_2 FILLER_0_134_744 ();
 sg13g2_fill_1 FILLER_0_134_746 ();
 sg13g2_fill_2 FILLER_0_134_752 ();
 sg13g2_fill_4 FILLER_0_134_759 ();
 sg13g2_fill_1 FILLER_0_134_763 ();
 sg13g2_fill_8 FILLER_0_134_768 ();
 sg13g2_fill_2 FILLER_0_134_776 ();
 sg13g2_fill_1 FILLER_0_134_778 ();
 sg13g2_fill_8 FILLER_0_134_784 ();
 sg13g2_fill_2 FILLER_0_134_792 ();
 sg13g2_fill_8 FILLER_0_134_820 ();
 sg13g2_fill_1 FILLER_0_134_828 ();
 sg13g2_fill_2 FILLER_0_134_839 ();
 sg13g2_fill_4 FILLER_0_134_849 ();
 sg13g2_fill_1 FILLER_0_134_853 ();
 sg13g2_fill_8 FILLER_0_134_862 ();
 sg13g2_fill_8 FILLER_0_134_876 ();
 sg13g2_fill_8 FILLER_0_134_884 ();
 sg13g2_fill_4 FILLER_0_134_892 ();
 sg13g2_fill_8 FILLER_0_134_901 ();
 sg13g2_fill_4 FILLER_0_134_909 ();
 sg13g2_fill_2 FILLER_0_134_917 ();
 sg13g2_fill_4 FILLER_0_134_924 ();
 sg13g2_fill_2 FILLER_0_134_928 ();
 sg13g2_fill_1 FILLER_0_134_930 ();
 sg13g2_fill_8 FILLER_0_134_941 ();
 sg13g2_fill_8 FILLER_0_134_949 ();
 sg13g2_fill_8 FILLER_0_134_957 ();
 sg13g2_fill_8 FILLER_0_134_965 ();
 sg13g2_fill_8 FILLER_0_134_973 ();
 sg13g2_fill_8 FILLER_0_134_981 ();
 sg13g2_fill_4 FILLER_0_134_989 ();
 sg13g2_fill_2 FILLER_0_134_993 ();
 sg13g2_fill_4 FILLER_0_134_1000 ();
 sg13g2_fill_4 FILLER_0_134_1008 ();
 sg13g2_fill_1 FILLER_0_134_1012 ();
 sg13g2_fill_8 FILLER_0_134_1020 ();
 sg13g2_fill_4 FILLER_0_134_1028 ();
 sg13g2_fill_2 FILLER_0_134_1032 ();
 sg13g2_fill_1 FILLER_0_134_1034 ();
 sg13g2_fill_2 FILLER_0_134_1041 ();
 sg13g2_fill_4 FILLER_0_134_1047 ();
 sg13g2_fill_2 FILLER_0_134_1058 ();
 sg13g2_fill_2 FILLER_0_134_1067 ();
 sg13g2_fill_4 FILLER_0_134_1095 ();
 sg13g2_fill_2 FILLER_0_134_1099 ();
 sg13g2_fill_8 FILLER_0_134_1106 ();
 sg13g2_fill_2 FILLER_0_134_1114 ();
 sg13g2_fill_1 FILLER_0_134_1116 ();
 sg13g2_fill_2 FILLER_0_134_1123 ();
 sg13g2_fill_8 FILLER_0_134_1130 ();
 sg13g2_fill_2 FILLER_0_134_1138 ();
 sg13g2_fill_2 FILLER_0_134_1145 ();
 sg13g2_fill_8 FILLER_0_134_1173 ();
 sg13g2_fill_8 FILLER_0_134_1181 ();
 sg13g2_fill_2 FILLER_0_134_1189 ();
 sg13g2_fill_1 FILLER_0_134_1191 ();
 sg13g2_fill_2 FILLER_0_134_1200 ();
 sg13g2_fill_8 FILLER_0_134_1207 ();
 sg13g2_fill_8 FILLER_0_134_1223 ();
 sg13g2_fill_1 FILLER_0_134_1231 ();
 sg13g2_fill_8 FILLER_0_134_1242 ();
 sg13g2_fill_8 FILLER_0_134_1250 ();
 sg13g2_fill_4 FILLER_0_134_1258 ();
 sg13g2_fill_2 FILLER_0_134_1262 ();
 sg13g2_fill_2 FILLER_0_134_1272 ();
 sg13g2_fill_4 FILLER_0_134_1278 ();
 sg13g2_fill_4 FILLER_0_134_1290 ();
 sg13g2_fill_2 FILLER_0_134_1294 ();
 sg13g2_fill_1 FILLER_0_134_1296 ();
 sg13g2_fill_8 FILLER_0_135_0 ();
 sg13g2_fill_8 FILLER_0_135_8 ();
 sg13g2_fill_8 FILLER_0_135_16 ();
 sg13g2_fill_8 FILLER_0_135_24 ();
 sg13g2_fill_8 FILLER_0_135_32 ();
 sg13g2_fill_8 FILLER_0_135_40 ();
 sg13g2_fill_8 FILLER_0_135_48 ();
 sg13g2_fill_8 FILLER_0_135_56 ();
 sg13g2_fill_8 FILLER_0_135_64 ();
 sg13g2_fill_8 FILLER_0_135_72 ();
 sg13g2_fill_8 FILLER_0_135_80 ();
 sg13g2_fill_8 FILLER_0_135_88 ();
 sg13g2_fill_8 FILLER_0_135_96 ();
 sg13g2_fill_8 FILLER_0_135_104 ();
 sg13g2_fill_8 FILLER_0_135_112 ();
 sg13g2_fill_8 FILLER_0_135_120 ();
 sg13g2_fill_8 FILLER_0_135_128 ();
 sg13g2_fill_8 FILLER_0_135_136 ();
 sg13g2_fill_8 FILLER_0_135_144 ();
 sg13g2_fill_8 FILLER_0_135_152 ();
 sg13g2_fill_8 FILLER_0_135_160 ();
 sg13g2_fill_8 FILLER_0_135_168 ();
 sg13g2_fill_8 FILLER_0_135_176 ();
 sg13g2_fill_8 FILLER_0_135_184 ();
 sg13g2_fill_8 FILLER_0_135_192 ();
 sg13g2_fill_8 FILLER_0_135_200 ();
 sg13g2_fill_8 FILLER_0_135_208 ();
 sg13g2_fill_8 FILLER_0_135_216 ();
 sg13g2_fill_8 FILLER_0_135_224 ();
 sg13g2_fill_8 FILLER_0_135_232 ();
 sg13g2_fill_8 FILLER_0_135_240 ();
 sg13g2_fill_8 FILLER_0_135_248 ();
 sg13g2_fill_8 FILLER_0_135_256 ();
 sg13g2_fill_8 FILLER_0_135_264 ();
 sg13g2_fill_8 FILLER_0_135_272 ();
 sg13g2_fill_8 FILLER_0_135_280 ();
 sg13g2_fill_8 FILLER_0_135_288 ();
 sg13g2_fill_2 FILLER_0_135_296 ();
 sg13g2_fill_1 FILLER_0_135_298 ();
 sg13g2_fill_4 FILLER_0_135_325 ();
 sg13g2_fill_2 FILLER_0_135_329 ();
 sg13g2_fill_2 FILLER_0_135_335 ();
 sg13g2_fill_8 FILLER_0_135_358 ();
 sg13g2_fill_8 FILLER_0_135_366 ();
 sg13g2_fill_8 FILLER_0_135_374 ();
 sg13g2_fill_4 FILLER_0_135_382 ();
 sg13g2_fill_2 FILLER_0_135_386 ();
 sg13g2_fill_1 FILLER_0_135_388 ();
 sg13g2_fill_4 FILLER_0_135_399 ();
 sg13g2_fill_4 FILLER_0_135_408 ();
 sg13g2_fill_4 FILLER_0_135_416 ();
 sg13g2_fill_4 FILLER_0_135_428 ();
 sg13g2_fill_2 FILLER_0_135_432 ();
 sg13g2_fill_2 FILLER_0_135_438 ();
 sg13g2_fill_4 FILLER_0_135_466 ();
 sg13g2_fill_2 FILLER_0_135_470 ();
 sg13g2_fill_1 FILLER_0_135_472 ();
 sg13g2_fill_4 FILLER_0_135_499 ();
 sg13g2_fill_1 FILLER_0_135_503 ();
 sg13g2_fill_8 FILLER_0_135_511 ();
 sg13g2_fill_8 FILLER_0_135_519 ();
 sg13g2_fill_4 FILLER_0_135_527 ();
 sg13g2_fill_2 FILLER_0_135_531 ();
 sg13g2_fill_8 FILLER_0_135_537 ();
 sg13g2_fill_8 FILLER_0_135_545 ();
 sg13g2_fill_4 FILLER_0_135_553 ();
 sg13g2_fill_1 FILLER_0_135_557 ();
 sg13g2_fill_8 FILLER_0_135_584 ();
 sg13g2_fill_8 FILLER_0_135_592 ();
 sg13g2_fill_8 FILLER_0_135_600 ();
 sg13g2_fill_8 FILLER_0_135_608 ();
 sg13g2_fill_2 FILLER_0_135_616 ();
 sg13g2_fill_1 FILLER_0_135_618 ();
 sg13g2_fill_8 FILLER_0_135_645 ();
 sg13g2_fill_4 FILLER_0_135_653 ();
 sg13g2_fill_2 FILLER_0_135_657 ();
 sg13g2_fill_1 FILLER_0_135_659 ();
 sg13g2_fill_4 FILLER_0_135_665 ();
 sg13g2_fill_2 FILLER_0_135_675 ();
 sg13g2_fill_1 FILLER_0_135_677 ();
 sg13g2_fill_4 FILLER_0_135_683 ();
 sg13g2_fill_4 FILLER_0_135_693 ();
 sg13g2_fill_2 FILLER_0_135_697 ();
 sg13g2_fill_8 FILLER_0_135_720 ();
 sg13g2_fill_8 FILLER_0_135_728 ();
 sg13g2_fill_8 FILLER_0_135_736 ();
 sg13g2_fill_8 FILLER_0_135_744 ();
 sg13g2_fill_4 FILLER_0_135_757 ();
 sg13g2_fill_2 FILLER_0_135_761 ();
 sg13g2_fill_8 FILLER_0_135_789 ();
 sg13g2_fill_8 FILLER_0_135_797 ();
 sg13g2_fill_4 FILLER_0_135_805 ();
 sg13g2_fill_1 FILLER_0_135_809 ();
 sg13g2_fill_8 FILLER_0_135_815 ();
 sg13g2_fill_8 FILLER_0_135_823 ();
 sg13g2_fill_2 FILLER_0_135_831 ();
 sg13g2_fill_2 FILLER_0_135_837 ();
 sg13g2_fill_1 FILLER_0_135_839 ();
 sg13g2_fill_8 FILLER_0_135_846 ();
 sg13g2_fill_4 FILLER_0_135_854 ();
 sg13g2_fill_1 FILLER_0_135_858 ();
 sg13g2_fill_2 FILLER_0_135_864 ();
 sg13g2_fill_1 FILLER_0_135_866 ();
 sg13g2_fill_8 FILLER_0_135_871 ();
 sg13g2_fill_8 FILLER_0_135_879 ();
 sg13g2_fill_8 FILLER_0_135_887 ();
 sg13g2_fill_8 FILLER_0_135_895 ();
 sg13g2_fill_8 FILLER_0_135_903 ();
 sg13g2_fill_2 FILLER_0_135_911 ();
 sg13g2_fill_1 FILLER_0_135_913 ();
 sg13g2_fill_4 FILLER_0_135_918 ();
 sg13g2_fill_4 FILLER_0_135_948 ();
 sg13g2_fill_2 FILLER_0_135_952 ();
 sg13g2_fill_1 FILLER_0_135_954 ();
 sg13g2_fill_8 FILLER_0_135_976 ();
 sg13g2_fill_8 FILLER_0_135_984 ();
 sg13g2_fill_1 FILLER_0_135_992 ();
 sg13g2_fill_8 FILLER_0_135_1019 ();
 sg13g2_fill_8 FILLER_0_135_1027 ();
 sg13g2_fill_8 FILLER_0_135_1035 ();
 sg13g2_fill_8 FILLER_0_135_1043 ();
 sg13g2_fill_4 FILLER_0_135_1051 ();
 sg13g2_fill_2 FILLER_0_135_1055 ();
 sg13g2_fill_1 FILLER_0_135_1057 ();
 sg13g2_fill_2 FILLER_0_135_1064 ();
 sg13g2_fill_1 FILLER_0_135_1066 ();
 sg13g2_fill_8 FILLER_0_135_1073 ();
 sg13g2_fill_2 FILLER_0_135_1081 ();
 sg13g2_fill_1 FILLER_0_135_1083 ();
 sg13g2_fill_2 FILLER_0_135_1090 ();
 sg13g2_fill_2 FILLER_0_135_1097 ();
 sg13g2_fill_2 FILLER_0_135_1125 ();
 sg13g2_fill_2 FILLER_0_135_1131 ();
 sg13g2_fill_1 FILLER_0_135_1133 ();
 sg13g2_fill_2 FILLER_0_135_1139 ();
 sg13g2_fill_8 FILLER_0_135_1167 ();
 sg13g2_fill_1 FILLER_0_135_1175 ();
 sg13g2_fill_8 FILLER_0_135_1181 ();
 sg13g2_fill_4 FILLER_0_135_1189 ();
 sg13g2_fill_1 FILLER_0_135_1193 ();
 sg13g2_fill_8 FILLER_0_135_1202 ();
 sg13g2_fill_8 FILLER_0_135_1210 ();
 sg13g2_fill_8 FILLER_0_135_1218 ();
 sg13g2_fill_4 FILLER_0_135_1226 ();
 sg13g2_fill_2 FILLER_0_135_1240 ();
 sg13g2_fill_2 FILLER_0_135_1268 ();
 sg13g2_fill_1 FILLER_0_135_1296 ();
 sg13g2_fill_8 FILLER_0_136_0 ();
 sg13g2_fill_8 FILLER_0_136_8 ();
 sg13g2_fill_8 FILLER_0_136_16 ();
 sg13g2_fill_8 FILLER_0_136_24 ();
 sg13g2_fill_8 FILLER_0_136_32 ();
 sg13g2_fill_8 FILLER_0_136_40 ();
 sg13g2_fill_8 FILLER_0_136_48 ();
 sg13g2_fill_8 FILLER_0_136_56 ();
 sg13g2_fill_8 FILLER_0_136_64 ();
 sg13g2_fill_8 FILLER_0_136_72 ();
 sg13g2_fill_8 FILLER_0_136_80 ();
 sg13g2_fill_8 FILLER_0_136_88 ();
 sg13g2_fill_8 FILLER_0_136_96 ();
 sg13g2_fill_8 FILLER_0_136_104 ();
 sg13g2_fill_8 FILLER_0_136_112 ();
 sg13g2_fill_8 FILLER_0_136_120 ();
 sg13g2_fill_8 FILLER_0_136_128 ();
 sg13g2_fill_8 FILLER_0_136_136 ();
 sg13g2_fill_8 FILLER_0_136_144 ();
 sg13g2_fill_8 FILLER_0_136_152 ();
 sg13g2_fill_8 FILLER_0_136_160 ();
 sg13g2_fill_8 FILLER_0_136_168 ();
 sg13g2_fill_8 FILLER_0_136_176 ();
 sg13g2_fill_8 FILLER_0_136_184 ();
 sg13g2_fill_8 FILLER_0_136_192 ();
 sg13g2_fill_8 FILLER_0_136_200 ();
 sg13g2_fill_8 FILLER_0_136_208 ();
 sg13g2_fill_8 FILLER_0_136_216 ();
 sg13g2_fill_8 FILLER_0_136_224 ();
 sg13g2_fill_8 FILLER_0_136_232 ();
 sg13g2_fill_8 FILLER_0_136_240 ();
 sg13g2_fill_8 FILLER_0_136_248 ();
 sg13g2_fill_8 FILLER_0_136_256 ();
 sg13g2_fill_8 FILLER_0_136_264 ();
 sg13g2_fill_8 FILLER_0_136_272 ();
 sg13g2_fill_8 FILLER_0_136_280 ();
 sg13g2_fill_2 FILLER_0_136_288 ();
 sg13g2_fill_1 FILLER_0_136_290 ();
 sg13g2_fill_4 FILLER_0_136_317 ();
 sg13g2_fill_2 FILLER_0_136_321 ();
 sg13g2_fill_8 FILLER_0_136_349 ();
 sg13g2_fill_8 FILLER_0_136_357 ();
 sg13g2_fill_8 FILLER_0_136_365 ();
 sg13g2_fill_8 FILLER_0_136_378 ();
 sg13g2_fill_8 FILLER_0_136_386 ();
 sg13g2_fill_8 FILLER_0_136_394 ();
 sg13g2_fill_8 FILLER_0_136_402 ();
 sg13g2_fill_2 FILLER_0_136_410 ();
 sg13g2_fill_1 FILLER_0_136_412 ();
 sg13g2_fill_2 FILLER_0_136_423 ();
 sg13g2_fill_4 FILLER_0_136_431 ();
 sg13g2_fill_8 FILLER_0_136_440 ();
 sg13g2_fill_8 FILLER_0_136_453 ();
 sg13g2_fill_8 FILLER_0_136_461 ();
 sg13g2_fill_8 FILLER_0_136_469 ();
 sg13g2_fill_8 FILLER_0_136_477 ();
 sg13g2_fill_8 FILLER_0_136_485 ();
 sg13g2_fill_8 FILLER_0_136_493 ();
 sg13g2_fill_2 FILLER_0_136_501 ();
 sg13g2_fill_4 FILLER_0_136_507 ();
 sg13g2_fill_1 FILLER_0_136_511 ();
 sg13g2_fill_2 FILLER_0_136_518 ();
 sg13g2_fill_1 FILLER_0_136_520 ();
 sg13g2_fill_4 FILLER_0_136_526 ();
 sg13g2_fill_2 FILLER_0_136_535 ();
 sg13g2_fill_8 FILLER_0_136_563 ();
 sg13g2_fill_8 FILLER_0_136_571 ();
 sg13g2_fill_4 FILLER_0_136_579 ();
 sg13g2_fill_4 FILLER_0_136_588 ();
 sg13g2_fill_1 FILLER_0_136_592 ();
 sg13g2_fill_8 FILLER_0_136_598 ();
 sg13g2_fill_8 FILLER_0_136_606 ();
 sg13g2_fill_2 FILLER_0_136_614 ();
 sg13g2_fill_1 FILLER_0_136_616 ();
 sg13g2_fill_8 FILLER_0_136_622 ();
 sg13g2_fill_8 FILLER_0_136_630 ();
 sg13g2_fill_8 FILLER_0_136_638 ();
 sg13g2_fill_8 FILLER_0_136_646 ();
 sg13g2_fill_8 FILLER_0_136_654 ();
 sg13g2_fill_2 FILLER_0_136_662 ();
 sg13g2_fill_2 FILLER_0_136_690 ();
 sg13g2_fill_2 FILLER_0_136_700 ();
 sg13g2_fill_2 FILLER_0_136_708 ();
 sg13g2_fill_8 FILLER_0_136_714 ();
 sg13g2_fill_8 FILLER_0_136_722 ();
 sg13g2_fill_8 FILLER_0_136_730 ();
 sg13g2_fill_2 FILLER_0_136_738 ();
 sg13g2_fill_1 FILLER_0_136_740 ();
 sg13g2_fill_2 FILLER_0_136_747 ();
 sg13g2_fill_8 FILLER_0_136_754 ();
 sg13g2_fill_8 FILLER_0_136_762 ();
 sg13g2_fill_1 FILLER_0_136_770 ();
 sg13g2_fill_2 FILLER_0_136_776 ();
 sg13g2_fill_8 FILLER_0_136_782 ();
 sg13g2_fill_8 FILLER_0_136_790 ();
 sg13g2_fill_8 FILLER_0_136_798 ();
 sg13g2_fill_8 FILLER_0_136_806 ();
 sg13g2_fill_8 FILLER_0_136_814 ();
 sg13g2_fill_2 FILLER_0_136_822 ();
 sg13g2_fill_2 FILLER_0_136_831 ();
 sg13g2_fill_8 FILLER_0_136_838 ();
 sg13g2_fill_4 FILLER_0_136_846 ();
 sg13g2_fill_2 FILLER_0_136_850 ();
 sg13g2_fill_2 FILLER_0_136_878 ();
 sg13g2_fill_8 FILLER_0_136_885 ();
 sg13g2_fill_8 FILLER_0_136_893 ();
 sg13g2_fill_8 FILLER_0_136_901 ();
 sg13g2_fill_2 FILLER_0_136_914 ();
 sg13g2_fill_1 FILLER_0_136_916 ();
 sg13g2_fill_2 FILLER_0_136_921 ();
 sg13g2_fill_8 FILLER_0_136_928 ();
 sg13g2_fill_4 FILLER_0_136_936 ();
 sg13g2_fill_2 FILLER_0_136_940 ();
 sg13g2_fill_1 FILLER_0_136_942 ();
 sg13g2_fill_2 FILLER_0_136_948 ();
 sg13g2_fill_2 FILLER_0_136_954 ();
 sg13g2_fill_2 FILLER_0_136_961 ();
 sg13g2_fill_4 FILLER_0_136_989 ();
 sg13g2_fill_2 FILLER_0_136_993 ();
 sg13g2_fill_1 FILLER_0_136_995 ();
 sg13g2_fill_8 FILLER_0_136_1001 ();
 sg13g2_fill_4 FILLER_0_136_1009 ();
 sg13g2_fill_2 FILLER_0_136_1013 ();
 sg13g2_fill_4 FILLER_0_136_1023 ();
 sg13g2_fill_8 FILLER_0_136_1031 ();
 sg13g2_fill_1 FILLER_0_136_1039 ();
 sg13g2_fill_4 FILLER_0_136_1045 ();
 sg13g2_fill_8 FILLER_0_136_1057 ();
 sg13g2_fill_8 FILLER_0_136_1065 ();
 sg13g2_fill_8 FILLER_0_136_1073 ();
 sg13g2_fill_8 FILLER_0_136_1081 ();
 sg13g2_fill_8 FILLER_0_136_1089 ();
 sg13g2_fill_2 FILLER_0_136_1097 ();
 sg13g2_fill_1 FILLER_0_136_1099 ();
 sg13g2_fill_2 FILLER_0_136_1105 ();
 sg13g2_fill_8 FILLER_0_136_1111 ();
 sg13g2_fill_4 FILLER_0_136_1119 ();
 sg13g2_fill_8 FILLER_0_136_1127 ();
 sg13g2_fill_8 FILLER_0_136_1135 ();
 sg13g2_fill_8 FILLER_0_136_1143 ();
 sg13g2_fill_8 FILLER_0_136_1151 ();
 sg13g2_fill_2 FILLER_0_136_1159 ();
 sg13g2_fill_1 FILLER_0_136_1161 ();
 sg13g2_fill_8 FILLER_0_136_1183 ();
 sg13g2_fill_8 FILLER_0_136_1191 ();
 sg13g2_fill_8 FILLER_0_136_1199 ();
 sg13g2_fill_8 FILLER_0_136_1207 ();
 sg13g2_fill_8 FILLER_0_136_1215 ();
 sg13g2_fill_8 FILLER_0_136_1223 ();
 sg13g2_fill_8 FILLER_0_136_1231 ();
 sg13g2_fill_8 FILLER_0_136_1239 ();
 sg13g2_fill_8 FILLER_0_136_1247 ();
 sg13g2_fill_2 FILLER_0_136_1255 ();
 sg13g2_fill_2 FILLER_0_136_1267 ();
 sg13g2_fill_8 FILLER_0_136_1279 ();
 sg13g2_fill_8 FILLER_0_136_1287 ();
 sg13g2_fill_2 FILLER_0_136_1295 ();
 sg13g2_fill_8 FILLER_0_137_0 ();
 sg13g2_fill_8 FILLER_0_137_8 ();
 sg13g2_fill_8 FILLER_0_137_16 ();
 sg13g2_fill_8 FILLER_0_137_24 ();
 sg13g2_fill_8 FILLER_0_137_32 ();
 sg13g2_fill_8 FILLER_0_137_40 ();
 sg13g2_fill_8 FILLER_0_137_48 ();
 sg13g2_fill_8 FILLER_0_137_56 ();
 sg13g2_fill_8 FILLER_0_137_64 ();
 sg13g2_fill_8 FILLER_0_137_72 ();
 sg13g2_fill_8 FILLER_0_137_80 ();
 sg13g2_fill_8 FILLER_0_137_88 ();
 sg13g2_fill_8 FILLER_0_137_96 ();
 sg13g2_fill_8 FILLER_0_137_104 ();
 sg13g2_fill_8 FILLER_0_137_112 ();
 sg13g2_fill_8 FILLER_0_137_120 ();
 sg13g2_fill_8 FILLER_0_137_128 ();
 sg13g2_fill_8 FILLER_0_137_136 ();
 sg13g2_fill_8 FILLER_0_137_144 ();
 sg13g2_fill_8 FILLER_0_137_152 ();
 sg13g2_fill_8 FILLER_0_137_160 ();
 sg13g2_fill_8 FILLER_0_137_168 ();
 sg13g2_fill_8 FILLER_0_137_176 ();
 sg13g2_fill_8 FILLER_0_137_184 ();
 sg13g2_fill_8 FILLER_0_137_192 ();
 sg13g2_fill_8 FILLER_0_137_200 ();
 sg13g2_fill_8 FILLER_0_137_208 ();
 sg13g2_fill_8 FILLER_0_137_216 ();
 sg13g2_fill_8 FILLER_0_137_224 ();
 sg13g2_fill_8 FILLER_0_137_232 ();
 sg13g2_fill_8 FILLER_0_137_240 ();
 sg13g2_fill_8 FILLER_0_137_248 ();
 sg13g2_fill_8 FILLER_0_137_256 ();
 sg13g2_fill_8 FILLER_0_137_264 ();
 sg13g2_fill_8 FILLER_0_137_272 ();
 sg13g2_fill_8 FILLER_0_137_280 ();
 sg13g2_fill_4 FILLER_0_137_288 ();
 sg13g2_fill_2 FILLER_0_137_292 ();
 sg13g2_fill_2 FILLER_0_137_299 ();
 sg13g2_fill_8 FILLER_0_137_305 ();
 sg13g2_fill_2 FILLER_0_137_313 ();
 sg13g2_fill_1 FILLER_0_137_315 ();
 sg13g2_fill_2 FILLER_0_137_322 ();
 sg13g2_fill_2 FILLER_0_137_329 ();
 sg13g2_fill_1 FILLER_0_137_331 ();
 sg13g2_fill_2 FILLER_0_137_353 ();
 sg13g2_fill_8 FILLER_0_137_360 ();
 sg13g2_fill_8 FILLER_0_137_368 ();
 sg13g2_fill_2 FILLER_0_137_380 ();
 sg13g2_fill_2 FILLER_0_137_387 ();
 sg13g2_fill_8 FILLER_0_137_393 ();
 sg13g2_fill_4 FILLER_0_137_401 ();
 sg13g2_fill_1 FILLER_0_137_405 ();
 sg13g2_fill_4 FILLER_0_137_418 ();
 sg13g2_fill_1 FILLER_0_137_422 ();
 sg13g2_fill_2 FILLER_0_137_428 ();
 sg13g2_fill_2 FILLER_0_137_434 ();
 sg13g2_fill_2 FILLER_0_137_440 ();
 sg13g2_fill_1 FILLER_0_137_442 ();
 sg13g2_fill_2 FILLER_0_137_448 ();
 sg13g2_fill_2 FILLER_0_137_455 ();
 sg13g2_fill_4 FILLER_0_137_462 ();
 sg13g2_fill_2 FILLER_0_137_466 ();
 sg13g2_fill_8 FILLER_0_137_494 ();
 sg13g2_fill_4 FILLER_0_137_508 ();
 sg13g2_fill_2 FILLER_0_137_512 ();
 sg13g2_fill_1 FILLER_0_137_514 ();
 sg13g2_fill_8 FILLER_0_137_520 ();
 sg13g2_fill_8 FILLER_0_137_528 ();
 sg13g2_fill_8 FILLER_0_137_536 ();
 sg13g2_fill_8 FILLER_0_137_544 ();
 sg13g2_fill_4 FILLER_0_137_552 ();
 sg13g2_fill_1 FILLER_0_137_556 ();
 sg13g2_fill_8 FILLER_0_137_567 ();
 sg13g2_fill_4 FILLER_0_137_579 ();
 sg13g2_fill_2 FILLER_0_137_583 ();
 sg13g2_fill_4 FILLER_0_137_590 ();
 sg13g2_fill_8 FILLER_0_137_599 ();
 sg13g2_fill_8 FILLER_0_137_607 ();
 sg13g2_fill_8 FILLER_0_137_615 ();
 sg13g2_fill_4 FILLER_0_137_623 ();
 sg13g2_fill_2 FILLER_0_137_633 ();
 sg13g2_fill_8 FILLER_0_137_640 ();
 sg13g2_fill_8 FILLER_0_137_648 ();
 sg13g2_fill_2 FILLER_0_137_660 ();
 sg13g2_fill_2 FILLER_0_137_667 ();
 sg13g2_fill_2 FILLER_0_137_673 ();
 sg13g2_fill_8 FILLER_0_137_680 ();
 sg13g2_fill_1 FILLER_0_137_688 ();
 sg13g2_fill_2 FILLER_0_137_697 ();
 sg13g2_fill_4 FILLER_0_137_707 ();
 sg13g2_fill_2 FILLER_0_137_711 ();
 sg13g2_fill_4 FILLER_0_137_718 ();
 sg13g2_fill_2 FILLER_0_137_722 ();
 sg13g2_fill_1 FILLER_0_137_724 ();
 sg13g2_fill_8 FILLER_0_137_751 ();
 sg13g2_fill_8 FILLER_0_137_759 ();
 sg13g2_fill_8 FILLER_0_137_767 ();
 sg13g2_fill_8 FILLER_0_137_775 ();
 sg13g2_fill_8 FILLER_0_137_783 ();
 sg13g2_fill_8 FILLER_0_137_791 ();
 sg13g2_fill_8 FILLER_0_137_799 ();
 sg13g2_fill_8 FILLER_0_137_813 ();
 sg13g2_fill_4 FILLER_0_137_821 ();
 sg13g2_fill_2 FILLER_0_137_825 ();
 sg13g2_fill_8 FILLER_0_137_853 ();
 sg13g2_fill_8 FILLER_0_137_861 ();
 sg13g2_fill_2 FILLER_0_137_874 ();
 sg13g2_fill_8 FILLER_0_137_880 ();
 sg13g2_fill_8 FILLER_0_137_888 ();
 sg13g2_fill_8 FILLER_0_137_896 ();
 sg13g2_fill_8 FILLER_0_137_904 ();
 sg13g2_fill_4 FILLER_0_137_912 ();
 sg13g2_fill_1 FILLER_0_137_916 ();
 sg13g2_fill_8 FILLER_0_137_943 ();
 sg13g2_fill_8 FILLER_0_137_951 ();
 sg13g2_fill_8 FILLER_0_137_959 ();
 sg13g2_fill_8 FILLER_0_137_967 ();
 sg13g2_fill_8 FILLER_0_137_975 ();
 sg13g2_fill_2 FILLER_0_137_983 ();
 sg13g2_fill_2 FILLER_0_137_995 ();
 sg13g2_fill_2 FILLER_0_137_1002 ();
 sg13g2_fill_8 FILLER_0_137_1009 ();
 sg13g2_fill_4 FILLER_0_137_1022 ();
 sg13g2_fill_2 FILLER_0_137_1026 ();
 sg13g2_fill_4 FILLER_0_137_1033 ();
 sg13g2_fill_2 FILLER_0_137_1042 ();
 sg13g2_fill_8 FILLER_0_137_1054 ();
 sg13g2_fill_8 FILLER_0_137_1062 ();
 sg13g2_fill_8 FILLER_0_137_1070 ();
 sg13g2_fill_8 FILLER_0_137_1078 ();
 sg13g2_fill_8 FILLER_0_137_1086 ();
 sg13g2_fill_8 FILLER_0_137_1094 ();
 sg13g2_fill_8 FILLER_0_137_1102 ();
 sg13g2_fill_8 FILLER_0_137_1110 ();
 sg13g2_fill_8 FILLER_0_137_1118 ();
 sg13g2_fill_8 FILLER_0_137_1126 ();
 sg13g2_fill_8 FILLER_0_137_1134 ();
 sg13g2_fill_8 FILLER_0_137_1142 ();
 sg13g2_fill_8 FILLER_0_137_1150 ();
 sg13g2_fill_8 FILLER_0_137_1158 ();
 sg13g2_fill_8 FILLER_0_137_1166 ();
 sg13g2_fill_8 FILLER_0_137_1174 ();
 sg13g2_fill_2 FILLER_0_137_1182 ();
 sg13g2_fill_2 FILLER_0_137_1210 ();
 sg13g2_fill_8 FILLER_0_137_1217 ();
 sg13g2_fill_8 FILLER_0_137_1225 ();
 sg13g2_fill_8 FILLER_0_137_1233 ();
 sg13g2_fill_8 FILLER_0_137_1241 ();
 sg13g2_fill_8 FILLER_0_137_1249 ();
 sg13g2_fill_8 FILLER_0_137_1257 ();
 sg13g2_fill_8 FILLER_0_137_1265 ();
 sg13g2_fill_8 FILLER_0_137_1273 ();
 sg13g2_fill_8 FILLER_0_137_1281 ();
 sg13g2_fill_8 FILLER_0_137_1289 ();
 sg13g2_fill_8 FILLER_0_138_0 ();
 sg13g2_fill_8 FILLER_0_138_8 ();
 sg13g2_fill_8 FILLER_0_138_16 ();
 sg13g2_fill_8 FILLER_0_138_24 ();
 sg13g2_fill_8 FILLER_0_138_32 ();
 sg13g2_fill_8 FILLER_0_138_40 ();
 sg13g2_fill_8 FILLER_0_138_48 ();
 sg13g2_fill_8 FILLER_0_138_56 ();
 sg13g2_fill_8 FILLER_0_138_64 ();
 sg13g2_fill_8 FILLER_0_138_72 ();
 sg13g2_fill_8 FILLER_0_138_80 ();
 sg13g2_fill_8 FILLER_0_138_88 ();
 sg13g2_fill_8 FILLER_0_138_96 ();
 sg13g2_fill_8 FILLER_0_138_104 ();
 sg13g2_fill_8 FILLER_0_138_112 ();
 sg13g2_fill_8 FILLER_0_138_120 ();
 sg13g2_fill_8 FILLER_0_138_128 ();
 sg13g2_fill_8 FILLER_0_138_136 ();
 sg13g2_fill_8 FILLER_0_138_144 ();
 sg13g2_fill_8 FILLER_0_138_152 ();
 sg13g2_fill_8 FILLER_0_138_160 ();
 sg13g2_fill_8 FILLER_0_138_168 ();
 sg13g2_fill_8 FILLER_0_138_176 ();
 sg13g2_fill_8 FILLER_0_138_184 ();
 sg13g2_fill_8 FILLER_0_138_192 ();
 sg13g2_fill_8 FILLER_0_138_200 ();
 sg13g2_fill_8 FILLER_0_138_208 ();
 sg13g2_fill_8 FILLER_0_138_216 ();
 sg13g2_fill_8 FILLER_0_138_224 ();
 sg13g2_fill_8 FILLER_0_138_232 ();
 sg13g2_fill_8 FILLER_0_138_240 ();
 sg13g2_fill_8 FILLER_0_138_248 ();
 sg13g2_fill_8 FILLER_0_138_256 ();
 sg13g2_fill_8 FILLER_0_138_264 ();
 sg13g2_fill_8 FILLER_0_138_272 ();
 sg13g2_fill_8 FILLER_0_138_280 ();
 sg13g2_fill_8 FILLER_0_138_288 ();
 sg13g2_fill_8 FILLER_0_138_296 ();
 sg13g2_fill_8 FILLER_0_138_304 ();
 sg13g2_fill_8 FILLER_0_138_312 ();
 sg13g2_fill_8 FILLER_0_138_320 ();
 sg13g2_fill_8 FILLER_0_138_328 ();
 sg13g2_fill_8 FILLER_0_138_336 ();
 sg13g2_fill_8 FILLER_0_138_344 ();
 sg13g2_fill_8 FILLER_0_138_352 ();
 sg13g2_fill_4 FILLER_0_138_360 ();
 sg13g2_fill_2 FILLER_0_138_390 ();
 sg13g2_fill_8 FILLER_0_138_397 ();
 sg13g2_fill_1 FILLER_0_138_405 ();
 sg13g2_fill_2 FILLER_0_138_410 ();
 sg13g2_fill_2 FILLER_0_138_417 ();
 sg13g2_fill_1 FILLER_0_138_419 ();
 sg13g2_fill_4 FILLER_0_138_425 ();
 sg13g2_fill_2 FILLER_0_138_429 ();
 sg13g2_fill_4 FILLER_0_138_434 ();
 sg13g2_fill_1 FILLER_0_138_438 ();
 sg13g2_fill_2 FILLER_0_138_445 ();
 sg13g2_fill_2 FILLER_0_138_454 ();
 sg13g2_fill_1 FILLER_0_138_456 ();
 sg13g2_fill_4 FILLER_0_138_465 ();
 sg13g2_fill_2 FILLER_0_138_469 ();
 sg13g2_fill_1 FILLER_0_138_471 ();
 sg13g2_fill_4 FILLER_0_138_498 ();
 sg13g2_fill_8 FILLER_0_138_507 ();
 sg13g2_fill_2 FILLER_0_138_515 ();
 sg13g2_fill_1 FILLER_0_138_517 ();
 sg13g2_fill_8 FILLER_0_138_523 ();
 sg13g2_fill_8 FILLER_0_138_531 ();
 sg13g2_fill_8 FILLER_0_138_539 ();
 sg13g2_fill_8 FILLER_0_138_547 ();
 sg13g2_fill_8 FILLER_0_138_555 ();
 sg13g2_fill_8 FILLER_0_138_563 ();
 sg13g2_fill_8 FILLER_0_138_571 ();
 sg13g2_fill_8 FILLER_0_138_579 ();
 sg13g2_fill_4 FILLER_0_138_587 ();
 sg13g2_fill_8 FILLER_0_138_598 ();
 sg13g2_fill_4 FILLER_0_138_606 ();
 sg13g2_fill_2 FILLER_0_138_610 ();
 sg13g2_fill_2 FILLER_0_138_638 ();
 sg13g2_fill_4 FILLER_0_138_644 ();
 sg13g2_fill_2 FILLER_0_138_648 ();
 sg13g2_fill_2 FILLER_0_138_655 ();
 sg13g2_fill_8 FILLER_0_138_661 ();
 sg13g2_fill_2 FILLER_0_138_669 ();
 sg13g2_fill_1 FILLER_0_138_671 ();
 sg13g2_fill_2 FILLER_0_138_677 ();
 sg13g2_fill_8 FILLER_0_138_684 ();
 sg13g2_fill_2 FILLER_0_138_692 ();
 sg13g2_fill_1 FILLER_0_138_694 ();
 sg13g2_fill_8 FILLER_0_138_700 ();
 sg13g2_fill_8 FILLER_0_138_708 ();
 sg13g2_fill_8 FILLER_0_138_716 ();
 sg13g2_fill_4 FILLER_0_138_724 ();
 sg13g2_fill_2 FILLER_0_138_733 ();
 sg13g2_fill_2 FILLER_0_138_739 ();
 sg13g2_fill_8 FILLER_0_138_746 ();
 sg13g2_fill_2 FILLER_0_138_754 ();
 sg13g2_fill_1 FILLER_0_138_756 ();
 sg13g2_fill_2 FILLER_0_138_762 ();
 sg13g2_fill_8 FILLER_0_138_770 ();
 sg13g2_fill_8 FILLER_0_138_778 ();
 sg13g2_fill_4 FILLER_0_138_786 ();
 sg13g2_fill_2 FILLER_0_138_790 ();
 sg13g2_fill_1 FILLER_0_138_792 ();
 sg13g2_fill_8 FILLER_0_138_799 ();
 sg13g2_fill_8 FILLER_0_138_807 ();
 sg13g2_fill_8 FILLER_0_138_815 ();
 sg13g2_fill_2 FILLER_0_138_823 ();
 sg13g2_fill_1 FILLER_0_138_825 ();
 sg13g2_fill_8 FILLER_0_138_832 ();
 sg13g2_fill_8 FILLER_0_138_840 ();
 sg13g2_fill_8 FILLER_0_138_848 ();
 sg13g2_fill_2 FILLER_0_138_861 ();
 sg13g2_fill_4 FILLER_0_138_889 ();
 sg13g2_fill_1 FILLER_0_138_893 ();
 sg13g2_fill_2 FILLER_0_138_898 ();
 sg13g2_fill_2 FILLER_0_138_926 ();
 sg13g2_fill_2 FILLER_0_138_933 ();
 sg13g2_fill_8 FILLER_0_138_939 ();
 sg13g2_fill_1 FILLER_0_138_947 ();
 sg13g2_fill_2 FILLER_0_138_953 ();
 sg13g2_fill_2 FILLER_0_138_981 ();
 sg13g2_fill_8 FILLER_0_138_1004 ();
 sg13g2_fill_4 FILLER_0_138_1012 ();
 sg13g2_fill_2 FILLER_0_138_1042 ();
 sg13g2_fill_2 FILLER_0_138_1049 ();
 sg13g2_fill_4 FILLER_0_138_1055 ();
 sg13g2_fill_2 FILLER_0_138_1064 ();
 sg13g2_fill_8 FILLER_0_138_1092 ();
 sg13g2_fill_4 FILLER_0_138_1100 ();
 sg13g2_fill_1 FILLER_0_138_1104 ();
 sg13g2_fill_2 FILLER_0_138_1110 ();
 sg13g2_fill_4 FILLER_0_138_1116 ();
 sg13g2_fill_1 FILLER_0_138_1120 ();
 sg13g2_fill_4 FILLER_0_138_1126 ();
 sg13g2_fill_2 FILLER_0_138_1130 ();
 sg13g2_fill_1 FILLER_0_138_1132 ();
 sg13g2_fill_2 FILLER_0_138_1138 ();
 sg13g2_fill_8 FILLER_0_138_1166 ();
 sg13g2_fill_4 FILLER_0_138_1174 ();
 sg13g2_fill_1 FILLER_0_138_1178 ();
 sg13g2_fill_4 FILLER_0_138_1183 ();
 sg13g2_fill_8 FILLER_0_138_1213 ();
 sg13g2_fill_8 FILLER_0_138_1221 ();
 sg13g2_fill_8 FILLER_0_138_1229 ();
 sg13g2_fill_8 FILLER_0_138_1237 ();
 sg13g2_fill_8 FILLER_0_138_1245 ();
 sg13g2_fill_8 FILLER_0_138_1253 ();
 sg13g2_fill_8 FILLER_0_138_1261 ();
 sg13g2_fill_8 FILLER_0_138_1269 ();
 sg13g2_fill_8 FILLER_0_138_1277 ();
 sg13g2_fill_8 FILLER_0_138_1285 ();
 sg13g2_fill_4 FILLER_0_138_1293 ();
 sg13g2_fill_8 FILLER_0_139_0 ();
 sg13g2_fill_8 FILLER_0_139_8 ();
 sg13g2_fill_8 FILLER_0_139_16 ();
 sg13g2_fill_8 FILLER_0_139_24 ();
 sg13g2_fill_8 FILLER_0_139_32 ();
 sg13g2_fill_8 FILLER_0_139_40 ();
 sg13g2_fill_8 FILLER_0_139_48 ();
 sg13g2_fill_8 FILLER_0_139_56 ();
 sg13g2_fill_8 FILLER_0_139_64 ();
 sg13g2_fill_8 FILLER_0_139_72 ();
 sg13g2_fill_8 FILLER_0_139_80 ();
 sg13g2_fill_8 FILLER_0_139_88 ();
 sg13g2_fill_8 FILLER_0_139_96 ();
 sg13g2_fill_8 FILLER_0_139_104 ();
 sg13g2_fill_8 FILLER_0_139_112 ();
 sg13g2_fill_8 FILLER_0_139_120 ();
 sg13g2_fill_8 FILLER_0_139_128 ();
 sg13g2_fill_8 FILLER_0_139_136 ();
 sg13g2_fill_8 FILLER_0_139_144 ();
 sg13g2_fill_8 FILLER_0_139_152 ();
 sg13g2_fill_8 FILLER_0_139_160 ();
 sg13g2_fill_8 FILLER_0_139_168 ();
 sg13g2_fill_8 FILLER_0_139_176 ();
 sg13g2_fill_8 FILLER_0_139_184 ();
 sg13g2_fill_8 FILLER_0_139_192 ();
 sg13g2_fill_8 FILLER_0_139_200 ();
 sg13g2_fill_8 FILLER_0_139_208 ();
 sg13g2_fill_8 FILLER_0_139_216 ();
 sg13g2_fill_8 FILLER_0_139_224 ();
 sg13g2_fill_8 FILLER_0_139_232 ();
 sg13g2_fill_8 FILLER_0_139_240 ();
 sg13g2_fill_8 FILLER_0_139_248 ();
 sg13g2_fill_8 FILLER_0_139_256 ();
 sg13g2_fill_8 FILLER_0_139_264 ();
 sg13g2_fill_8 FILLER_0_139_272 ();
 sg13g2_fill_8 FILLER_0_139_280 ();
 sg13g2_fill_8 FILLER_0_139_288 ();
 sg13g2_fill_4 FILLER_0_139_296 ();
 sg13g2_fill_1 FILLER_0_139_300 ();
 sg13g2_fill_2 FILLER_0_139_306 ();
 sg13g2_fill_8 FILLER_0_139_312 ();
 sg13g2_fill_8 FILLER_0_139_320 ();
 sg13g2_fill_1 FILLER_0_139_328 ();
 sg13g2_fill_8 FILLER_0_139_337 ();
 sg13g2_fill_2 FILLER_0_139_371 ();
 sg13g2_fill_8 FILLER_0_139_377 ();
 sg13g2_fill_4 FILLER_0_139_385 ();
 sg13g2_fill_2 FILLER_0_139_389 ();
 sg13g2_fill_1 FILLER_0_139_391 ();
 sg13g2_fill_2 FILLER_0_139_396 ();
 sg13g2_fill_4 FILLER_0_139_403 ();
 sg13g2_fill_2 FILLER_0_139_407 ();
 sg13g2_fill_8 FILLER_0_139_417 ();
 sg13g2_fill_8 FILLER_0_139_425 ();
 sg13g2_fill_8 FILLER_0_139_433 ();
 sg13g2_fill_4 FILLER_0_139_441 ();
 sg13g2_fill_2 FILLER_0_139_445 ();
 sg13g2_fill_1 FILLER_0_139_447 ();
 sg13g2_fill_8 FILLER_0_139_453 ();
 sg13g2_fill_8 FILLER_0_139_461 ();
 sg13g2_fill_2 FILLER_0_139_474 ();
 sg13g2_fill_2 FILLER_0_139_480 ();
 sg13g2_fill_1 FILLER_0_139_482 ();
 sg13g2_fill_8 FILLER_0_139_487 ();
 sg13g2_fill_8 FILLER_0_139_495 ();
 sg13g2_fill_4 FILLER_0_139_503 ();
 sg13g2_fill_2 FILLER_0_139_507 ();
 sg13g2_fill_1 FILLER_0_139_509 ();
 sg13g2_fill_2 FILLER_0_139_536 ();
 sg13g2_fill_4 FILLER_0_139_564 ();
 sg13g2_fill_2 FILLER_0_139_568 ();
 sg13g2_fill_1 FILLER_0_139_570 ();
 sg13g2_fill_8 FILLER_0_139_597 ();
 sg13g2_fill_2 FILLER_0_139_610 ();
 sg13g2_fill_4 FILLER_0_139_616 ();
 sg13g2_fill_2 FILLER_0_139_620 ();
 sg13g2_fill_8 FILLER_0_139_627 ();
 sg13g2_fill_8 FILLER_0_139_635 ();
 sg13g2_fill_4 FILLER_0_139_643 ();
 sg13g2_fill_8 FILLER_0_139_673 ();
 sg13g2_fill_8 FILLER_0_139_707 ();
 sg13g2_fill_4 FILLER_0_139_715 ();
 sg13g2_fill_2 FILLER_0_139_719 ();
 sg13g2_fill_2 FILLER_0_139_747 ();
 sg13g2_fill_2 FILLER_0_139_753 ();
 sg13g2_fill_4 FILLER_0_139_760 ();
 sg13g2_fill_2 FILLER_0_139_764 ();
 sg13g2_fill_4 FILLER_0_139_772 ();
 sg13g2_fill_4 FILLER_0_139_781 ();
 sg13g2_fill_2 FILLER_0_139_785 ();
 sg13g2_fill_1 FILLER_0_139_787 ();
 sg13g2_fill_8 FILLER_0_139_814 ();
 sg13g2_fill_8 FILLER_0_139_822 ();
 sg13g2_fill_4 FILLER_0_139_830 ();
 sg13g2_fill_2 FILLER_0_139_838 ();
 sg13g2_fill_4 FILLER_0_139_845 ();
 sg13g2_fill_2 FILLER_0_139_849 ();
 sg13g2_fill_1 FILLER_0_139_851 ();
 sg13g2_fill_8 FILLER_0_139_857 ();
 sg13g2_fill_8 FILLER_0_139_865 ();
 sg13g2_fill_8 FILLER_0_139_873 ();
 sg13g2_fill_1 FILLER_0_139_881 ();
 sg13g2_fill_8 FILLER_0_139_887 ();
 sg13g2_fill_4 FILLER_0_139_895 ();
 sg13g2_fill_1 FILLER_0_139_899 ();
 sg13g2_fill_4 FILLER_0_139_905 ();
 sg13g2_fill_1 FILLER_0_139_909 ();
 sg13g2_fill_8 FILLER_0_139_920 ();
 sg13g2_fill_8 FILLER_0_139_928 ();
 sg13g2_fill_8 FILLER_0_139_936 ();
 sg13g2_fill_8 FILLER_0_139_944 ();
 sg13g2_fill_4 FILLER_0_139_952 ();
 sg13g2_fill_1 FILLER_0_139_956 ();
 sg13g2_fill_2 FILLER_0_139_962 ();
 sg13g2_fill_8 FILLER_0_139_968 ();
 sg13g2_fill_4 FILLER_0_139_976 ();
 sg13g2_fill_2 FILLER_0_139_980 ();
 sg13g2_fill_1 FILLER_0_139_982 ();
 sg13g2_fill_8 FILLER_0_139_993 ();
 sg13g2_fill_8 FILLER_0_139_1001 ();
 sg13g2_fill_4 FILLER_0_139_1009 ();
 sg13g2_fill_1 FILLER_0_139_1013 ();
 sg13g2_fill_2 FILLER_0_139_1019 ();
 sg13g2_fill_1 FILLER_0_139_1021 ();
 sg13g2_fill_8 FILLER_0_139_1027 ();
 sg13g2_fill_8 FILLER_0_139_1035 ();
 sg13g2_fill_8 FILLER_0_139_1043 ();
 sg13g2_fill_4 FILLER_0_139_1051 ();
 sg13g2_fill_1 FILLER_0_139_1055 ();
 sg13g2_fill_4 FILLER_0_139_1061 ();
 sg13g2_fill_4 FILLER_0_139_1073 ();
 sg13g2_fill_2 FILLER_0_139_1077 ();
 sg13g2_fill_1 FILLER_0_139_1079 ();
 sg13g2_fill_8 FILLER_0_139_1085 ();
 sg13g2_fill_8 FILLER_0_139_1093 ();
 sg13g2_fill_2 FILLER_0_139_1101 ();
 sg13g2_fill_2 FILLER_0_139_1129 ();
 sg13g2_fill_2 FILLER_0_139_1135 ();
 sg13g2_fill_8 FILLER_0_139_1142 ();
 sg13g2_fill_8 FILLER_0_139_1150 ();
 sg13g2_fill_8 FILLER_0_139_1158 ();
 sg13g2_fill_8 FILLER_0_139_1166 ();
 sg13g2_fill_2 FILLER_0_139_1178 ();
 sg13g2_fill_2 FILLER_0_139_1185 ();
 sg13g2_fill_2 FILLER_0_139_1208 ();
 sg13g2_fill_4 FILLER_0_139_1214 ();
 sg13g2_fill_2 FILLER_0_139_1223 ();
 sg13g2_fill_2 FILLER_0_139_1251 ();
 sg13g2_fill_8 FILLER_0_139_1257 ();
 sg13g2_fill_8 FILLER_0_139_1265 ();
 sg13g2_fill_8 FILLER_0_139_1273 ();
 sg13g2_fill_8 FILLER_0_139_1281 ();
 sg13g2_fill_8 FILLER_0_139_1289 ();
 sg13g2_fill_8 FILLER_0_140_0 ();
 sg13g2_fill_8 FILLER_0_140_8 ();
 sg13g2_fill_8 FILLER_0_140_16 ();
 sg13g2_fill_8 FILLER_0_140_24 ();
 sg13g2_fill_8 FILLER_0_140_32 ();
 sg13g2_fill_8 FILLER_0_140_40 ();
 sg13g2_fill_8 FILLER_0_140_48 ();
 sg13g2_fill_8 FILLER_0_140_56 ();
 sg13g2_fill_8 FILLER_0_140_64 ();
 sg13g2_fill_8 FILLER_0_140_72 ();
 sg13g2_fill_8 FILLER_0_140_80 ();
 sg13g2_fill_8 FILLER_0_140_88 ();
 sg13g2_fill_8 FILLER_0_140_96 ();
 sg13g2_fill_8 FILLER_0_140_104 ();
 sg13g2_fill_8 FILLER_0_140_112 ();
 sg13g2_fill_8 FILLER_0_140_120 ();
 sg13g2_fill_8 FILLER_0_140_128 ();
 sg13g2_fill_8 FILLER_0_140_136 ();
 sg13g2_fill_8 FILLER_0_140_144 ();
 sg13g2_fill_8 FILLER_0_140_152 ();
 sg13g2_fill_8 FILLER_0_140_160 ();
 sg13g2_fill_8 FILLER_0_140_168 ();
 sg13g2_fill_8 FILLER_0_140_176 ();
 sg13g2_fill_8 FILLER_0_140_184 ();
 sg13g2_fill_8 FILLER_0_140_192 ();
 sg13g2_fill_8 FILLER_0_140_200 ();
 sg13g2_fill_8 FILLER_0_140_208 ();
 sg13g2_fill_8 FILLER_0_140_216 ();
 sg13g2_fill_8 FILLER_0_140_224 ();
 sg13g2_fill_8 FILLER_0_140_232 ();
 sg13g2_fill_8 FILLER_0_140_240 ();
 sg13g2_fill_8 FILLER_0_140_248 ();
 sg13g2_fill_8 FILLER_0_140_256 ();
 sg13g2_fill_8 FILLER_0_140_264 ();
 sg13g2_fill_8 FILLER_0_140_272 ();
 sg13g2_fill_8 FILLER_0_140_280 ();
 sg13g2_fill_2 FILLER_0_140_288 ();
 sg13g2_fill_1 FILLER_0_140_290 ();
 sg13g2_fill_2 FILLER_0_140_317 ();
 sg13g2_fill_2 FILLER_0_140_324 ();
 sg13g2_fill_1 FILLER_0_140_326 ();
 sg13g2_fill_2 FILLER_0_140_333 ();
 sg13g2_fill_4 FILLER_0_140_356 ();
 sg13g2_fill_2 FILLER_0_140_360 ();
 sg13g2_fill_1 FILLER_0_140_362 ();
 sg13g2_fill_2 FILLER_0_140_371 ();
 sg13g2_fill_1 FILLER_0_140_373 ();
 sg13g2_fill_2 FILLER_0_140_395 ();
 sg13g2_fill_4 FILLER_0_140_423 ();
 sg13g2_fill_2 FILLER_0_140_432 ();
 sg13g2_fill_8 FILLER_0_140_438 ();
 sg13g2_fill_8 FILLER_0_140_451 ();
 sg13g2_fill_8 FILLER_0_140_459 ();
 sg13g2_fill_8 FILLER_0_140_467 ();
 sg13g2_fill_4 FILLER_0_140_475 ();
 sg13g2_fill_1 FILLER_0_140_479 ();
 sg13g2_fill_8 FILLER_0_140_485 ();
 sg13g2_fill_8 FILLER_0_140_493 ();
 sg13g2_fill_8 FILLER_0_140_501 ();
 sg13g2_fill_2 FILLER_0_140_513 ();
 sg13g2_fill_1 FILLER_0_140_515 ();
 sg13g2_fill_2 FILLER_0_140_521 ();
 sg13g2_fill_1 FILLER_0_140_523 ();
 sg13g2_fill_2 FILLER_0_140_528 ();
 sg13g2_fill_1 FILLER_0_140_530 ();
 sg13g2_fill_4 FILLER_0_140_535 ();
 sg13g2_fill_2 FILLER_0_140_560 ();
 sg13g2_fill_4 FILLER_0_140_566 ();
 sg13g2_fill_1 FILLER_0_140_570 ();
 sg13g2_fill_4 FILLER_0_140_576 ();
 sg13g2_fill_2 FILLER_0_140_580 ();
 sg13g2_fill_1 FILLER_0_140_582 ();
 sg13g2_fill_4 FILLER_0_140_587 ();
 sg13g2_fill_2 FILLER_0_140_591 ();
 sg13g2_fill_1 FILLER_0_140_593 ();
 sg13g2_fill_4 FILLER_0_140_598 ();
 sg13g2_fill_1 FILLER_0_140_602 ();
 sg13g2_fill_4 FILLER_0_140_629 ();
 sg13g2_fill_1 FILLER_0_140_633 ();
 sg13g2_fill_4 FILLER_0_140_655 ();
 sg13g2_fill_8 FILLER_0_140_666 ();
 sg13g2_fill_4 FILLER_0_140_674 ();
 sg13g2_fill_1 FILLER_0_140_678 ();
 sg13g2_fill_8 FILLER_0_140_683 ();
 sg13g2_fill_2 FILLER_0_140_691 ();
 sg13g2_fill_1 FILLER_0_140_693 ();
 sg13g2_fill_2 FILLER_0_140_700 ();
 sg13g2_fill_8 FILLER_0_140_707 ();
 sg13g2_fill_8 FILLER_0_140_715 ();
 sg13g2_fill_8 FILLER_0_140_723 ();
 sg13g2_fill_1 FILLER_0_140_731 ();
 sg13g2_fill_2 FILLER_0_140_737 ();
 sg13g2_fill_8 FILLER_0_140_743 ();
 sg13g2_fill_8 FILLER_0_140_751 ();
 sg13g2_fill_4 FILLER_0_140_759 ();
 sg13g2_fill_2 FILLER_0_140_763 ();
 sg13g2_fill_8 FILLER_0_140_771 ();
 sg13g2_fill_2 FILLER_0_140_779 ();
 sg13g2_fill_1 FILLER_0_140_781 ();
 sg13g2_fill_2 FILLER_0_140_787 ();
 sg13g2_fill_1 FILLER_0_140_789 ();
 sg13g2_fill_2 FILLER_0_140_795 ();
 sg13g2_fill_2 FILLER_0_140_802 ();
 sg13g2_fill_8 FILLER_0_140_808 ();
 sg13g2_fill_8 FILLER_0_140_816 ();
 sg13g2_fill_8 FILLER_0_140_824 ();
 sg13g2_fill_8 FILLER_0_140_832 ();
 sg13g2_fill_8 FILLER_0_140_840 ();
 sg13g2_fill_4 FILLER_0_140_848 ();
 sg13g2_fill_1 FILLER_0_140_852 ();
 sg13g2_fill_4 FILLER_0_140_859 ();
 sg13g2_fill_2 FILLER_0_140_863 ();
 sg13g2_fill_1 FILLER_0_140_865 ();
 sg13g2_fill_4 FILLER_0_140_874 ();
 sg13g2_fill_1 FILLER_0_140_878 ();
 sg13g2_fill_2 FILLER_0_140_885 ();
 sg13g2_fill_4 FILLER_0_140_913 ();
 sg13g2_fill_2 FILLER_0_140_917 ();
 sg13g2_fill_8 FILLER_0_140_924 ();
 sg13g2_fill_8 FILLER_0_140_942 ();
 sg13g2_fill_8 FILLER_0_140_950 ();
 sg13g2_fill_1 FILLER_0_140_958 ();
 sg13g2_fill_4 FILLER_0_140_964 ();
 sg13g2_fill_2 FILLER_0_140_968 ();
 sg13g2_fill_2 FILLER_0_140_980 ();
 sg13g2_fill_1 FILLER_0_140_982 ();
 sg13g2_fill_4 FILLER_0_140_1009 ();
 sg13g2_fill_4 FILLER_0_140_1023 ();
 sg13g2_fill_1 FILLER_0_140_1027 ();
 sg13g2_fill_2 FILLER_0_140_1033 ();
 sg13g2_fill_2 FILLER_0_140_1039 ();
 sg13g2_fill_2 FILLER_0_140_1046 ();
 sg13g2_fill_1 FILLER_0_140_1048 ();
 sg13g2_fill_2 FILLER_0_140_1055 ();
 sg13g2_fill_8 FILLER_0_140_1063 ();
 sg13g2_fill_2 FILLER_0_140_1071 ();
 sg13g2_fill_8 FILLER_0_140_1079 ();
 sg13g2_fill_8 FILLER_0_140_1087 ();
 sg13g2_fill_8 FILLER_0_140_1095 ();
 sg13g2_fill_8 FILLER_0_140_1103 ();
 sg13g2_fill_8 FILLER_0_140_1111 ();
 sg13g2_fill_8 FILLER_0_140_1119 ();
 sg13g2_fill_2 FILLER_0_140_1127 ();
 sg13g2_fill_8 FILLER_0_140_1139 ();
 sg13g2_fill_8 FILLER_0_140_1147 ();
 sg13g2_fill_8 FILLER_0_140_1155 ();
 sg13g2_fill_8 FILLER_0_140_1163 ();
 sg13g2_fill_2 FILLER_0_140_1171 ();
 sg13g2_fill_2 FILLER_0_140_1178 ();
 sg13g2_fill_2 FILLER_0_140_1206 ();
 sg13g2_fill_1 FILLER_0_140_1208 ();
 sg13g2_fill_2 FILLER_0_140_1214 ();
 sg13g2_fill_1 FILLER_0_140_1216 ();
 sg13g2_fill_2 FILLER_0_140_1222 ();
 sg13g2_fill_8 FILLER_0_140_1229 ();
 sg13g2_fill_1 FILLER_0_140_1237 ();
 sg13g2_fill_8 FILLER_0_140_1241 ();
 sg13g2_fill_2 FILLER_0_140_1249 ();
 sg13g2_fill_8 FILLER_0_140_1256 ();
 sg13g2_fill_8 FILLER_0_140_1264 ();
 sg13g2_fill_8 FILLER_0_140_1272 ();
 sg13g2_fill_8 FILLER_0_140_1280 ();
 sg13g2_fill_8 FILLER_0_140_1288 ();
 sg13g2_fill_1 FILLER_0_140_1296 ();
 sg13g2_fill_8 FILLER_0_141_0 ();
 sg13g2_fill_8 FILLER_0_141_8 ();
 sg13g2_fill_8 FILLER_0_141_16 ();
 sg13g2_fill_8 FILLER_0_141_24 ();
 sg13g2_fill_8 FILLER_0_141_32 ();
 sg13g2_fill_8 FILLER_0_141_40 ();
 sg13g2_fill_8 FILLER_0_141_48 ();
 sg13g2_fill_8 FILLER_0_141_56 ();
 sg13g2_fill_8 FILLER_0_141_64 ();
 sg13g2_fill_8 FILLER_0_141_72 ();
 sg13g2_fill_8 FILLER_0_141_80 ();
 sg13g2_fill_8 FILLER_0_141_88 ();
 sg13g2_fill_8 FILLER_0_141_96 ();
 sg13g2_fill_8 FILLER_0_141_104 ();
 sg13g2_fill_8 FILLER_0_141_112 ();
 sg13g2_fill_8 FILLER_0_141_120 ();
 sg13g2_fill_8 FILLER_0_141_128 ();
 sg13g2_fill_8 FILLER_0_141_136 ();
 sg13g2_fill_8 FILLER_0_141_144 ();
 sg13g2_fill_8 FILLER_0_141_152 ();
 sg13g2_fill_8 FILLER_0_141_160 ();
 sg13g2_fill_8 FILLER_0_141_168 ();
 sg13g2_fill_8 FILLER_0_141_176 ();
 sg13g2_fill_8 FILLER_0_141_184 ();
 sg13g2_fill_8 FILLER_0_141_192 ();
 sg13g2_fill_8 FILLER_0_141_200 ();
 sg13g2_fill_8 FILLER_0_141_208 ();
 sg13g2_fill_8 FILLER_0_141_216 ();
 sg13g2_fill_8 FILLER_0_141_224 ();
 sg13g2_fill_8 FILLER_0_141_232 ();
 sg13g2_fill_8 FILLER_0_141_240 ();
 sg13g2_fill_8 FILLER_0_141_248 ();
 sg13g2_fill_8 FILLER_0_141_256 ();
 sg13g2_fill_8 FILLER_0_141_264 ();
 sg13g2_fill_8 FILLER_0_141_272 ();
 sg13g2_fill_8 FILLER_0_141_280 ();
 sg13g2_fill_2 FILLER_0_141_292 ();
 sg13g2_fill_4 FILLER_0_141_299 ();
 sg13g2_fill_1 FILLER_0_141_303 ();
 sg13g2_fill_4 FILLER_0_141_330 ();
 sg13g2_fill_2 FILLER_0_141_334 ();
 sg13g2_fill_1 FILLER_0_141_336 ();
 sg13g2_fill_4 FILLER_0_141_341 ();
 sg13g2_fill_1 FILLER_0_141_345 ();
 sg13g2_fill_2 FILLER_0_141_350 ();
 sg13g2_fill_1 FILLER_0_141_352 ();
 sg13g2_fill_8 FILLER_0_141_379 ();
 sg13g2_fill_8 FILLER_0_141_387 ();
 sg13g2_fill_8 FILLER_0_141_395 ();
 sg13g2_fill_8 FILLER_0_141_403 ();
 sg13g2_fill_2 FILLER_0_141_411 ();
 sg13g2_fill_2 FILLER_0_141_417 ();
 sg13g2_fill_1 FILLER_0_141_419 ();
 sg13g2_fill_2 FILLER_0_141_424 ();
 sg13g2_fill_8 FILLER_0_141_452 ();
 sg13g2_fill_1 FILLER_0_141_460 ();
 sg13g2_fill_2 FILLER_0_141_487 ();
 sg13g2_fill_2 FILLER_0_141_510 ();
 sg13g2_fill_4 FILLER_0_141_517 ();
 sg13g2_fill_4 FILLER_0_141_525 ();
 sg13g2_fill_2 FILLER_0_141_529 ();
 sg13g2_fill_4 FILLER_0_141_536 ();
 sg13g2_fill_1 FILLER_0_141_540 ();
 sg13g2_fill_8 FILLER_0_141_545 ();
 sg13g2_fill_8 FILLER_0_141_553 ();
 sg13g2_fill_8 FILLER_0_141_561 ();
 sg13g2_fill_2 FILLER_0_141_574 ();
 sg13g2_fill_4 FILLER_0_141_584 ();
 sg13g2_fill_8 FILLER_0_141_596 ();
 sg13g2_fill_2 FILLER_0_141_610 ();
 sg13g2_fill_8 FILLER_0_141_617 ();
 sg13g2_fill_8 FILLER_0_141_625 ();
 sg13g2_fill_8 FILLER_0_141_633 ();
 sg13g2_fill_8 FILLER_0_141_641 ();
 sg13g2_fill_8 FILLER_0_141_649 ();
 sg13g2_fill_8 FILLER_0_141_657 ();
 sg13g2_fill_8 FILLER_0_141_665 ();
 sg13g2_fill_4 FILLER_0_141_673 ();
 sg13g2_fill_2 FILLER_0_141_681 ();
 sg13g2_fill_1 FILLER_0_141_683 ();
 sg13g2_fill_8 FILLER_0_141_710 ();
 sg13g2_fill_8 FILLER_0_141_718 ();
 sg13g2_fill_8 FILLER_0_141_726 ();
 sg13g2_fill_8 FILLER_0_141_734 ();
 sg13g2_fill_8 FILLER_0_141_742 ();
 sg13g2_fill_4 FILLER_0_141_750 ();
 sg13g2_fill_1 FILLER_0_141_754 ();
 sg13g2_fill_8 FILLER_0_141_760 ();
 sg13g2_fill_4 FILLER_0_141_768 ();
 sg13g2_fill_2 FILLER_0_141_772 ();
 sg13g2_fill_1 FILLER_0_141_774 ();
 sg13g2_fill_8 FILLER_0_141_780 ();
 sg13g2_fill_4 FILLER_0_141_788 ();
 sg13g2_fill_1 FILLER_0_141_792 ();
 sg13g2_fill_2 FILLER_0_141_798 ();
 sg13g2_fill_1 FILLER_0_141_800 ();
 sg13g2_fill_2 FILLER_0_141_805 ();
 sg13g2_fill_2 FILLER_0_141_833 ();
 sg13g2_fill_1 FILLER_0_141_835 ();
 sg13g2_fill_8 FILLER_0_141_862 ();
 sg13g2_fill_8 FILLER_0_141_870 ();
 sg13g2_fill_8 FILLER_0_141_878 ();
 sg13g2_fill_4 FILLER_0_141_886 ();
 sg13g2_fill_2 FILLER_0_141_890 ();
 sg13g2_fill_8 FILLER_0_141_896 ();
 sg13g2_fill_8 FILLER_0_141_904 ();
 sg13g2_fill_8 FILLER_0_141_912 ();
 sg13g2_fill_8 FILLER_0_141_925 ();
 sg13g2_fill_2 FILLER_0_141_954 ();
 sg13g2_fill_8 FILLER_0_141_982 ();
 sg13g2_fill_2 FILLER_0_141_995 ();
 sg13g2_fill_8 FILLER_0_141_1001 ();
 sg13g2_fill_8 FILLER_0_141_1009 ();
 sg13g2_fill_1 FILLER_0_141_1017 ();
 sg13g2_fill_2 FILLER_0_141_1044 ();
 sg13g2_fill_8 FILLER_0_141_1051 ();
 sg13g2_fill_8 FILLER_0_141_1059 ();
 sg13g2_fill_8 FILLER_0_141_1067 ();
 sg13g2_fill_8 FILLER_0_141_1080 ();
 sg13g2_fill_1 FILLER_0_141_1088 ();
 sg13g2_fill_4 FILLER_0_141_1093 ();
 sg13g2_fill_1 FILLER_0_141_1097 ();
 sg13g2_fill_8 FILLER_0_141_1102 ();
 sg13g2_fill_2 FILLER_0_141_1115 ();
 sg13g2_fill_2 FILLER_0_141_1143 ();
 sg13g2_fill_8 FILLER_0_141_1150 ();
 sg13g2_fill_4 FILLER_0_141_1158 ();
 sg13g2_fill_1 FILLER_0_141_1162 ();
 sg13g2_fill_8 FILLER_0_141_1189 ();
 sg13g2_fill_2 FILLER_0_141_1218 ();
 sg13g2_fill_8 FILLER_0_141_1225 ();
 sg13g2_fill_8 FILLER_0_141_1233 ();
 sg13g2_fill_8 FILLER_0_141_1241 ();
 sg13g2_fill_8 FILLER_0_141_1254 ();
 sg13g2_fill_8 FILLER_0_141_1262 ();
 sg13g2_fill_8 FILLER_0_141_1270 ();
 sg13g2_fill_8 FILLER_0_141_1278 ();
 sg13g2_fill_8 FILLER_0_141_1286 ();
 sg13g2_fill_2 FILLER_0_141_1294 ();
 sg13g2_fill_1 FILLER_0_141_1296 ();
 sg13g2_fill_8 FILLER_0_142_0 ();
 sg13g2_fill_8 FILLER_0_142_8 ();
 sg13g2_fill_8 FILLER_0_142_16 ();
 sg13g2_fill_8 FILLER_0_142_24 ();
 sg13g2_fill_8 FILLER_0_142_32 ();
 sg13g2_fill_8 FILLER_0_142_40 ();
 sg13g2_fill_8 FILLER_0_142_48 ();
 sg13g2_fill_8 FILLER_0_142_56 ();
 sg13g2_fill_8 FILLER_0_142_64 ();
 sg13g2_fill_8 FILLER_0_142_72 ();
 sg13g2_fill_8 FILLER_0_142_80 ();
 sg13g2_fill_8 FILLER_0_142_88 ();
 sg13g2_fill_8 FILLER_0_142_96 ();
 sg13g2_fill_8 FILLER_0_142_104 ();
 sg13g2_fill_8 FILLER_0_142_112 ();
 sg13g2_fill_8 FILLER_0_142_120 ();
 sg13g2_fill_8 FILLER_0_142_128 ();
 sg13g2_fill_8 FILLER_0_142_136 ();
 sg13g2_fill_8 FILLER_0_142_144 ();
 sg13g2_fill_8 FILLER_0_142_152 ();
 sg13g2_fill_8 FILLER_0_142_160 ();
 sg13g2_fill_8 FILLER_0_142_168 ();
 sg13g2_fill_8 FILLER_0_142_176 ();
 sg13g2_fill_8 FILLER_0_142_184 ();
 sg13g2_fill_8 FILLER_0_142_192 ();
 sg13g2_fill_8 FILLER_0_142_200 ();
 sg13g2_fill_8 FILLER_0_142_208 ();
 sg13g2_fill_8 FILLER_0_142_216 ();
 sg13g2_fill_8 FILLER_0_142_224 ();
 sg13g2_fill_8 FILLER_0_142_232 ();
 sg13g2_fill_8 FILLER_0_142_240 ();
 sg13g2_fill_8 FILLER_0_142_248 ();
 sg13g2_fill_8 FILLER_0_142_256 ();
 sg13g2_fill_8 FILLER_0_142_264 ();
 sg13g2_fill_8 FILLER_0_142_272 ();
 sg13g2_fill_8 FILLER_0_142_280 ();
 sg13g2_fill_8 FILLER_0_142_288 ();
 sg13g2_fill_4 FILLER_0_142_296 ();
 sg13g2_fill_2 FILLER_0_142_305 ();
 sg13g2_fill_1 FILLER_0_142_307 ();
 sg13g2_fill_4 FILLER_0_142_312 ();
 sg13g2_fill_1 FILLER_0_142_316 ();
 sg13g2_fill_4 FILLER_0_142_321 ();
 sg13g2_fill_1 FILLER_0_142_325 ();
 sg13g2_fill_2 FILLER_0_142_334 ();
 sg13g2_fill_4 FILLER_0_142_341 ();
 sg13g2_fill_8 FILLER_0_142_350 ();
 sg13g2_fill_8 FILLER_0_142_358 ();
 sg13g2_fill_8 FILLER_0_142_366 ();
 sg13g2_fill_2 FILLER_0_142_374 ();
 sg13g2_fill_2 FILLER_0_142_402 ();
 sg13g2_fill_4 FILLER_0_142_409 ();
 sg13g2_fill_1 FILLER_0_142_413 ();
 sg13g2_fill_8 FILLER_0_142_435 ();
 sg13g2_fill_8 FILLER_0_142_443 ();
 sg13g2_fill_8 FILLER_0_142_451 ();
 sg13g2_fill_2 FILLER_0_142_459 ();
 sg13g2_fill_1 FILLER_0_142_461 ();
 sg13g2_fill_4 FILLER_0_142_467 ();
 sg13g2_fill_1 FILLER_0_142_471 ();
 sg13g2_fill_2 FILLER_0_142_498 ();
 sg13g2_fill_8 FILLER_0_142_526 ();
 sg13g2_fill_8 FILLER_0_142_534 ();
 sg13g2_fill_8 FILLER_0_142_542 ();
 sg13g2_fill_8 FILLER_0_142_550 ();
 sg13g2_fill_8 FILLER_0_142_558 ();
 sg13g2_fill_8 FILLER_0_142_566 ();
 sg13g2_fill_8 FILLER_0_142_574 ();
 sg13g2_fill_8 FILLER_0_142_582 ();
 sg13g2_fill_8 FILLER_0_142_590 ();
 sg13g2_fill_8 FILLER_0_142_598 ();
 sg13g2_fill_8 FILLER_0_142_606 ();
 sg13g2_fill_8 FILLER_0_142_614 ();
 sg13g2_fill_8 FILLER_0_142_622 ();
 sg13g2_fill_8 FILLER_0_142_630 ();
 sg13g2_fill_8 FILLER_0_142_638 ();
 sg13g2_fill_8 FILLER_0_142_646 ();
 sg13g2_fill_8 FILLER_0_142_654 ();
 sg13g2_fill_2 FILLER_0_142_662 ();
 sg13g2_fill_8 FILLER_0_142_669 ();
 sg13g2_fill_8 FILLER_0_142_677 ();
 sg13g2_fill_2 FILLER_0_142_685 ();
 sg13g2_fill_1 FILLER_0_142_687 ();
 sg13g2_fill_8 FILLER_0_142_696 ();
 sg13g2_fill_8 FILLER_0_142_704 ();
 sg13g2_fill_8 FILLER_0_142_712 ();
 sg13g2_fill_2 FILLER_0_142_720 ();
 sg13g2_fill_1 FILLER_0_142_722 ();
 sg13g2_fill_2 FILLER_0_142_728 ();
 sg13g2_fill_1 FILLER_0_142_730 ();
 sg13g2_fill_2 FILLER_0_142_735 ();
 sg13g2_fill_1 FILLER_0_142_737 ();
 sg13g2_fill_2 FILLER_0_142_744 ();
 sg13g2_fill_1 FILLER_0_142_746 ();
 sg13g2_fill_8 FILLER_0_142_757 ();
 sg13g2_fill_4 FILLER_0_142_765 ();
 sg13g2_fill_2 FILLER_0_142_769 ();
 sg13g2_fill_1 FILLER_0_142_771 ();
 sg13g2_fill_4 FILLER_0_142_798 ();
 sg13g2_fill_2 FILLER_0_142_802 ();
 sg13g2_fill_8 FILLER_0_142_825 ();
 sg13g2_fill_4 FILLER_0_142_833 ();
 sg13g2_fill_2 FILLER_0_142_842 ();
 sg13g2_fill_1 FILLER_0_142_844 ();
 sg13g2_fill_8 FILLER_0_142_849 ();
 sg13g2_fill_8 FILLER_0_142_857 ();
 sg13g2_fill_8 FILLER_0_142_865 ();
 sg13g2_fill_8 FILLER_0_142_873 ();
 sg13g2_fill_8 FILLER_0_142_881 ();
 sg13g2_fill_8 FILLER_0_142_889 ();
 sg13g2_fill_4 FILLER_0_142_897 ();
 sg13g2_fill_2 FILLER_0_142_901 ();
 sg13g2_fill_1 FILLER_0_142_903 ();
 sg13g2_fill_4 FILLER_0_142_909 ();
 sg13g2_fill_2 FILLER_0_142_913 ();
 sg13g2_fill_1 FILLER_0_142_915 ();
 sg13g2_fill_2 FILLER_0_142_942 ();
 sg13g2_fill_4 FILLER_0_142_948 ();
 sg13g2_fill_2 FILLER_0_142_952 ();
 sg13g2_fill_1 FILLER_0_142_954 ();
 sg13g2_fill_8 FILLER_0_142_960 ();
 sg13g2_fill_8 FILLER_0_142_968 ();
 sg13g2_fill_8 FILLER_0_142_976 ();
 sg13g2_fill_8 FILLER_0_142_984 ();
 sg13g2_fill_8 FILLER_0_142_992 ();
 sg13g2_fill_8 FILLER_0_142_1005 ();
 sg13g2_fill_1 FILLER_0_142_1013 ();
 sg13g2_fill_8 FILLER_0_142_1018 ();
 sg13g2_fill_8 FILLER_0_142_1026 ();
 sg13g2_fill_8 FILLER_0_142_1034 ();
 sg13g2_fill_8 FILLER_0_142_1042 ();
 sg13g2_fill_8 FILLER_0_142_1050 ();
 sg13g2_fill_8 FILLER_0_142_1058 ();
 sg13g2_fill_8 FILLER_0_142_1066 ();
 sg13g2_fill_2 FILLER_0_142_1074 ();
 sg13g2_fill_1 FILLER_0_142_1076 ();
 sg13g2_fill_8 FILLER_0_142_1103 ();
 sg13g2_fill_2 FILLER_0_142_1111 ();
 sg13g2_fill_8 FILLER_0_142_1117 ();
 sg13g2_fill_8 FILLER_0_142_1125 ();
 sg13g2_fill_8 FILLER_0_142_1133 ();
 sg13g2_fill_2 FILLER_0_142_1141 ();
 sg13g2_fill_2 FILLER_0_142_1147 ();
 sg13g2_fill_1 FILLER_0_142_1149 ();
 sg13g2_fill_8 FILLER_0_142_1154 ();
 sg13g2_fill_4 FILLER_0_142_1162 ();
 sg13g2_fill_2 FILLER_0_142_1166 ();
 sg13g2_fill_1 FILLER_0_142_1168 ();
 sg13g2_fill_8 FILLER_0_142_1175 ();
 sg13g2_fill_8 FILLER_0_142_1183 ();
 sg13g2_fill_8 FILLER_0_142_1191 ();
 sg13g2_fill_1 FILLER_0_142_1199 ();
 sg13g2_fill_2 FILLER_0_142_1205 ();
 sg13g2_fill_8 FILLER_0_142_1212 ();
 sg13g2_fill_8 FILLER_0_142_1220 ();
 sg13g2_fill_8 FILLER_0_142_1228 ();
 sg13g2_fill_8 FILLER_0_142_1236 ();
 sg13g2_fill_8 FILLER_0_142_1244 ();
 sg13g2_fill_8 FILLER_0_142_1256 ();
 sg13g2_fill_8 FILLER_0_142_1264 ();
 sg13g2_fill_8 FILLER_0_142_1272 ();
 sg13g2_fill_8 FILLER_0_142_1280 ();
 sg13g2_fill_8 FILLER_0_142_1288 ();
 sg13g2_fill_1 FILLER_0_142_1296 ();
 sg13g2_fill_8 FILLER_0_143_0 ();
 sg13g2_fill_8 FILLER_0_143_8 ();
 sg13g2_fill_8 FILLER_0_143_16 ();
 sg13g2_fill_8 FILLER_0_143_24 ();
 sg13g2_fill_8 FILLER_0_143_32 ();
 sg13g2_fill_8 FILLER_0_143_40 ();
 sg13g2_fill_8 FILLER_0_143_48 ();
 sg13g2_fill_8 FILLER_0_143_56 ();
 sg13g2_fill_8 FILLER_0_143_64 ();
 sg13g2_fill_8 FILLER_0_143_72 ();
 sg13g2_fill_8 FILLER_0_143_80 ();
 sg13g2_fill_8 FILLER_0_143_88 ();
 sg13g2_fill_8 FILLER_0_143_96 ();
 sg13g2_fill_8 FILLER_0_143_104 ();
 sg13g2_fill_8 FILLER_0_143_112 ();
 sg13g2_fill_8 FILLER_0_143_120 ();
 sg13g2_fill_8 FILLER_0_143_128 ();
 sg13g2_fill_8 FILLER_0_143_136 ();
 sg13g2_fill_8 FILLER_0_143_144 ();
 sg13g2_fill_8 FILLER_0_143_152 ();
 sg13g2_fill_8 FILLER_0_143_160 ();
 sg13g2_fill_8 FILLER_0_143_168 ();
 sg13g2_fill_8 FILLER_0_143_176 ();
 sg13g2_fill_8 FILLER_0_143_184 ();
 sg13g2_fill_8 FILLER_0_143_192 ();
 sg13g2_fill_8 FILLER_0_143_200 ();
 sg13g2_fill_8 FILLER_0_143_208 ();
 sg13g2_fill_8 FILLER_0_143_216 ();
 sg13g2_fill_8 FILLER_0_143_224 ();
 sg13g2_fill_8 FILLER_0_143_232 ();
 sg13g2_fill_8 FILLER_0_143_240 ();
 sg13g2_fill_8 FILLER_0_143_248 ();
 sg13g2_fill_8 FILLER_0_143_256 ();
 sg13g2_fill_8 FILLER_0_143_264 ();
 sg13g2_fill_8 FILLER_0_143_272 ();
 sg13g2_fill_8 FILLER_0_143_280 ();
 sg13g2_fill_8 FILLER_0_143_288 ();
 sg13g2_fill_8 FILLER_0_143_296 ();
 sg13g2_fill_8 FILLER_0_143_304 ();
 sg13g2_fill_8 FILLER_0_143_312 ();
 sg13g2_fill_1 FILLER_0_143_320 ();
 sg13g2_fill_4 FILLER_0_143_326 ();
 sg13g2_fill_1 FILLER_0_143_330 ();
 sg13g2_fill_8 FILLER_0_143_336 ();
 sg13g2_fill_8 FILLER_0_143_344 ();
 sg13g2_fill_8 FILLER_0_143_352 ();
 sg13g2_fill_4 FILLER_0_143_360 ();
 sg13g2_fill_2 FILLER_0_143_364 ();
 sg13g2_fill_8 FILLER_0_143_370 ();
 sg13g2_fill_4 FILLER_0_143_378 ();
 sg13g2_fill_1 FILLER_0_143_382 ();
 sg13g2_fill_4 FILLER_0_143_388 ();
 sg13g2_fill_8 FILLER_0_143_396 ();
 sg13g2_fill_8 FILLER_0_143_404 ();
 sg13g2_fill_2 FILLER_0_143_412 ();
 sg13g2_fill_8 FILLER_0_143_440 ();
 sg13g2_fill_8 FILLER_0_143_448 ();
 sg13g2_fill_8 FILLER_0_143_456 ();
 sg13g2_fill_2 FILLER_0_143_464 ();
 sg13g2_fill_2 FILLER_0_143_470 ();
 sg13g2_fill_2 FILLER_0_143_477 ();
 sg13g2_fill_2 FILLER_0_143_483 ();
 sg13g2_fill_2 FILLER_0_143_506 ();
 sg13g2_fill_8 FILLER_0_143_513 ();
 sg13g2_fill_8 FILLER_0_143_521 ();
 sg13g2_fill_8 FILLER_0_143_529 ();
 sg13g2_fill_4 FILLER_0_143_542 ();
 sg13g2_fill_2 FILLER_0_143_546 ();
 sg13g2_fill_8 FILLER_0_143_574 ();
 sg13g2_fill_8 FILLER_0_143_582 ();
 sg13g2_fill_8 FILLER_0_143_590 ();
 sg13g2_fill_1 FILLER_0_143_598 ();
 sg13g2_fill_4 FILLER_0_143_625 ();
 sg13g2_fill_2 FILLER_0_143_629 ();
 sg13g2_fill_4 FILLER_0_143_637 ();
 sg13g2_fill_1 FILLER_0_143_641 ();
 sg13g2_fill_4 FILLER_0_143_668 ();
 sg13g2_fill_1 FILLER_0_143_672 ();
 sg13g2_fill_8 FILLER_0_143_678 ();
 sg13g2_fill_1 FILLER_0_143_686 ();
 sg13g2_fill_8 FILLER_0_143_692 ();
 sg13g2_fill_2 FILLER_0_143_700 ();
 sg13g2_fill_2 FILLER_0_143_706 ();
 sg13g2_fill_4 FILLER_0_143_713 ();
 sg13g2_fill_2 FILLER_0_143_717 ();
 sg13g2_fill_1 FILLER_0_143_719 ();
 sg13g2_fill_8 FILLER_0_143_746 ();
 sg13g2_fill_8 FILLER_0_143_758 ();
 sg13g2_fill_8 FILLER_0_143_766 ();
 sg13g2_fill_8 FILLER_0_143_774 ();
 sg13g2_fill_2 FILLER_0_143_808 ();
 sg13g2_fill_1 FILLER_0_143_810 ();
 sg13g2_fill_2 FILLER_0_143_816 ();
 sg13g2_fill_8 FILLER_0_143_822 ();
 sg13g2_fill_8 FILLER_0_143_830 ();
 sg13g2_fill_8 FILLER_0_143_838 ();
 sg13g2_fill_4 FILLER_0_143_846 ();
 sg13g2_fill_2 FILLER_0_143_850 ();
 sg13g2_fill_1 FILLER_0_143_852 ();
 sg13g2_fill_2 FILLER_0_143_863 ();
 sg13g2_fill_1 FILLER_0_143_865 ();
 sg13g2_fill_8 FILLER_0_143_872 ();
 sg13g2_fill_8 FILLER_0_143_880 ();
 sg13g2_fill_4 FILLER_0_143_888 ();
 sg13g2_fill_2 FILLER_0_143_892 ();
 sg13g2_fill_1 FILLER_0_143_894 ();
 sg13g2_fill_2 FILLER_0_143_921 ();
 sg13g2_fill_4 FILLER_0_143_927 ();
 sg13g2_fill_8 FILLER_0_143_935 ();
 sg13g2_fill_8 FILLER_0_143_943 ();
 sg13g2_fill_4 FILLER_0_143_951 ();
 sg13g2_fill_2 FILLER_0_143_955 ();
 sg13g2_fill_1 FILLER_0_143_957 ();
 sg13g2_fill_2 FILLER_0_143_963 ();
 sg13g2_fill_1 FILLER_0_143_965 ();
 sg13g2_fill_8 FILLER_0_143_971 ();
 sg13g2_fill_8 FILLER_0_143_979 ();
 sg13g2_fill_8 FILLER_0_143_987 ();
 sg13g2_fill_2 FILLER_0_143_995 ();
 sg13g2_fill_8 FILLER_0_143_1023 ();
 sg13g2_fill_2 FILLER_0_143_1031 ();
 sg13g2_fill_8 FILLER_0_143_1041 ();
 sg13g2_fill_8 FILLER_0_143_1049 ();
 sg13g2_fill_2 FILLER_0_143_1057 ();
 sg13g2_fill_1 FILLER_0_143_1059 ();
 sg13g2_fill_2 FILLER_0_143_1065 ();
 sg13g2_fill_2 FILLER_0_143_1071 ();
 sg13g2_fill_8 FILLER_0_143_1099 ();
 sg13g2_fill_8 FILLER_0_143_1107 ();
 sg13g2_fill_8 FILLER_0_143_1115 ();
 sg13g2_fill_8 FILLER_0_143_1123 ();
 sg13g2_fill_8 FILLER_0_143_1131 ();
 sg13g2_fill_4 FILLER_0_143_1139 ();
 sg13g2_fill_1 FILLER_0_143_1143 ();
 sg13g2_fill_8 FILLER_0_143_1154 ();
 sg13g2_fill_8 FILLER_0_143_1162 ();
 sg13g2_fill_2 FILLER_0_143_1170 ();
 sg13g2_fill_1 FILLER_0_143_1172 ();
 sg13g2_fill_2 FILLER_0_143_1179 ();
 sg13g2_fill_2 FILLER_0_143_1207 ();
 sg13g2_fill_4 FILLER_0_143_1214 ();
 sg13g2_fill_1 FILLER_0_143_1218 ();
 sg13g2_fill_8 FILLER_0_143_1223 ();
 sg13g2_fill_8 FILLER_0_143_1231 ();
 sg13g2_fill_4 FILLER_0_143_1239 ();
 sg13g2_fill_1 FILLER_0_143_1243 ();
 sg13g2_fill_8 FILLER_0_143_1270 ();
 sg13g2_fill_8 FILLER_0_143_1278 ();
 sg13g2_fill_8 FILLER_0_143_1286 ();
 sg13g2_fill_2 FILLER_0_143_1294 ();
 sg13g2_fill_1 FILLER_0_143_1296 ();
 sg13g2_fill_8 FILLER_0_144_0 ();
 sg13g2_fill_8 FILLER_0_144_8 ();
 sg13g2_fill_8 FILLER_0_144_16 ();
 sg13g2_fill_8 FILLER_0_144_24 ();
 sg13g2_fill_8 FILLER_0_144_32 ();
 sg13g2_fill_8 FILLER_0_144_40 ();
 sg13g2_fill_8 FILLER_0_144_48 ();
 sg13g2_fill_8 FILLER_0_144_56 ();
 sg13g2_fill_8 FILLER_0_144_64 ();
 sg13g2_fill_8 FILLER_0_144_72 ();
 sg13g2_fill_8 FILLER_0_144_80 ();
 sg13g2_fill_8 FILLER_0_144_88 ();
 sg13g2_fill_8 FILLER_0_144_96 ();
 sg13g2_fill_8 FILLER_0_144_104 ();
 sg13g2_fill_8 FILLER_0_144_112 ();
 sg13g2_fill_8 FILLER_0_144_120 ();
 sg13g2_fill_8 FILLER_0_144_128 ();
 sg13g2_fill_8 FILLER_0_144_136 ();
 sg13g2_fill_8 FILLER_0_144_144 ();
 sg13g2_fill_8 FILLER_0_144_152 ();
 sg13g2_fill_8 FILLER_0_144_160 ();
 sg13g2_fill_8 FILLER_0_144_168 ();
 sg13g2_fill_8 FILLER_0_144_176 ();
 sg13g2_fill_8 FILLER_0_144_184 ();
 sg13g2_fill_8 FILLER_0_144_192 ();
 sg13g2_fill_8 FILLER_0_144_200 ();
 sg13g2_fill_8 FILLER_0_144_208 ();
 sg13g2_fill_8 FILLER_0_144_216 ();
 sg13g2_fill_8 FILLER_0_144_224 ();
 sg13g2_fill_8 FILLER_0_144_232 ();
 sg13g2_fill_8 FILLER_0_144_240 ();
 sg13g2_fill_8 FILLER_0_144_248 ();
 sg13g2_fill_8 FILLER_0_144_256 ();
 sg13g2_fill_8 FILLER_0_144_264 ();
 sg13g2_fill_8 FILLER_0_144_272 ();
 sg13g2_fill_8 FILLER_0_144_280 ();
 sg13g2_fill_8 FILLER_0_144_288 ();
 sg13g2_fill_8 FILLER_0_144_296 ();
 sg13g2_fill_8 FILLER_0_144_304 ();
 sg13g2_fill_8 FILLER_0_144_312 ();
 sg13g2_fill_8 FILLER_0_144_320 ();
 sg13g2_fill_8 FILLER_0_144_328 ();
 sg13g2_fill_8 FILLER_0_144_336 ();
 sg13g2_fill_4 FILLER_0_144_344 ();
 sg13g2_fill_8 FILLER_0_144_352 ();
 sg13g2_fill_8 FILLER_0_144_360 ();
 sg13g2_fill_8 FILLER_0_144_368 ();
 sg13g2_fill_8 FILLER_0_144_376 ();
 sg13g2_fill_8 FILLER_0_144_384 ();
 sg13g2_fill_8 FILLER_0_144_392 ();
 sg13g2_fill_8 FILLER_0_144_400 ();
 sg13g2_fill_4 FILLER_0_144_408 ();
 sg13g2_fill_2 FILLER_0_144_417 ();
 sg13g2_fill_8 FILLER_0_144_423 ();
 sg13g2_fill_8 FILLER_0_144_431 ();
 sg13g2_fill_2 FILLER_0_144_439 ();
 sg13g2_fill_1 FILLER_0_144_441 ();
 sg13g2_fill_2 FILLER_0_144_448 ();
 sg13g2_fill_8 FILLER_0_144_458 ();
 sg13g2_fill_8 FILLER_0_144_466 ();
 sg13g2_fill_8 FILLER_0_144_474 ();
 sg13g2_fill_8 FILLER_0_144_482 ();
 sg13g2_fill_2 FILLER_0_144_490 ();
 sg13g2_fill_8 FILLER_0_144_497 ();
 sg13g2_fill_8 FILLER_0_144_505 ();
 sg13g2_fill_8 FILLER_0_144_513 ();
 sg13g2_fill_4 FILLER_0_144_521 ();
 sg13g2_fill_8 FILLER_0_144_530 ();
 sg13g2_fill_2 FILLER_0_144_542 ();
 sg13g2_fill_2 FILLER_0_144_548 ();
 sg13g2_fill_1 FILLER_0_144_550 ();
 sg13g2_fill_2 FILLER_0_144_572 ();
 sg13g2_fill_2 FILLER_0_144_579 ();
 sg13g2_fill_2 FILLER_0_144_585 ();
 sg13g2_fill_8 FILLER_0_144_591 ();
 sg13g2_fill_4 FILLER_0_144_599 ();
 sg13g2_fill_1 FILLER_0_144_603 ();
 sg13g2_fill_4 FILLER_0_144_609 ();
 sg13g2_fill_2 FILLER_0_144_639 ();
 sg13g2_fill_1 FILLER_0_144_641 ();
 sg13g2_fill_2 FILLER_0_144_647 ();
 sg13g2_fill_2 FILLER_0_144_670 ();
 sg13g2_fill_4 FILLER_0_144_698 ();
 sg13g2_fill_2 FILLER_0_144_702 ();
 sg13g2_fill_2 FILLER_0_144_730 ();
 sg13g2_fill_2 FILLER_0_144_736 ();
 sg13g2_fill_1 FILLER_0_144_738 ();
 sg13g2_fill_8 FILLER_0_144_743 ();
 sg13g2_fill_2 FILLER_0_144_751 ();
 sg13g2_fill_4 FILLER_0_144_758 ();
 sg13g2_fill_2 FILLER_0_144_762 ();
 sg13g2_fill_1 FILLER_0_144_764 ();
 sg13g2_fill_2 FILLER_0_144_771 ();
 sg13g2_fill_8 FILLER_0_144_777 ();
 sg13g2_fill_4 FILLER_0_144_785 ();
 sg13g2_fill_1 FILLER_0_144_789 ();
 sg13g2_fill_4 FILLER_0_144_795 ();
 sg13g2_fill_2 FILLER_0_144_799 ();
 sg13g2_fill_1 FILLER_0_144_801 ();
 sg13g2_fill_8 FILLER_0_144_806 ();
 sg13g2_fill_8 FILLER_0_144_814 ();
 sg13g2_fill_8 FILLER_0_144_827 ();
 sg13g2_fill_1 FILLER_0_144_835 ();
 sg13g2_fill_4 FILLER_0_144_857 ();
 sg13g2_fill_1 FILLER_0_144_861 ();
 sg13g2_fill_2 FILLER_0_144_866 ();
 sg13g2_fill_2 FILLER_0_144_872 ();
 sg13g2_fill_8 FILLER_0_144_879 ();
 sg13g2_fill_8 FILLER_0_144_887 ();
 sg13g2_fill_8 FILLER_0_144_895 ();
 sg13g2_fill_8 FILLER_0_144_903 ();
 sg13g2_fill_1 FILLER_0_144_911 ();
 sg13g2_fill_8 FILLER_0_144_938 ();
 sg13g2_fill_2 FILLER_0_144_946 ();
 sg13g2_fill_1 FILLER_0_144_948 ();
 sg13g2_fill_2 FILLER_0_144_954 ();
 sg13g2_fill_1 FILLER_0_144_956 ();
 sg13g2_fill_8 FILLER_0_144_961 ();
 sg13g2_fill_4 FILLER_0_144_969 ();
 sg13g2_fill_1 FILLER_0_144_973 ();
 sg13g2_fill_8 FILLER_0_144_981 ();
 sg13g2_fill_8 FILLER_0_144_989 ();
 sg13g2_fill_8 FILLER_0_144_997 ();
 sg13g2_fill_8 FILLER_0_144_1005 ();
 sg13g2_fill_4 FILLER_0_144_1013 ();
 sg13g2_fill_8 FILLER_0_144_1022 ();
 sg13g2_fill_8 FILLER_0_144_1030 ();
 sg13g2_fill_8 FILLER_0_144_1038 ();
 sg13g2_fill_2 FILLER_0_144_1046 ();
 sg13g2_fill_4 FILLER_0_144_1052 ();
 sg13g2_fill_8 FILLER_0_144_1062 ();
 sg13g2_fill_2 FILLER_0_144_1070 ();
 sg13g2_fill_1 FILLER_0_144_1072 ();
 sg13g2_fill_8 FILLER_0_144_1078 ();
 sg13g2_fill_1 FILLER_0_144_1086 ();
 sg13g2_fill_2 FILLER_0_144_1097 ();
 sg13g2_fill_8 FILLER_0_144_1109 ();
 sg13g2_fill_8 FILLER_0_144_1122 ();
 sg13g2_fill_2 FILLER_0_144_1130 ();
 sg13g2_fill_2 FILLER_0_144_1137 ();
 sg13g2_fill_4 FILLER_0_144_1143 ();
 sg13g2_fill_8 FILLER_0_144_1152 ();
 sg13g2_fill_8 FILLER_0_144_1160 ();
 sg13g2_fill_8 FILLER_0_144_1168 ();
 sg13g2_fill_2 FILLER_0_144_1176 ();
 sg13g2_fill_1 FILLER_0_144_1178 ();
 sg13g2_fill_2 FILLER_0_144_1184 ();
 sg13g2_fill_8 FILLER_0_144_1190 ();
 sg13g2_fill_4 FILLER_0_144_1198 ();
 sg13g2_fill_1 FILLER_0_144_1202 ();
 sg13g2_fill_8 FILLER_0_144_1224 ();
 sg13g2_fill_2 FILLER_0_144_1258 ();
 sg13g2_fill_8 FILLER_0_144_1265 ();
 sg13g2_fill_8 FILLER_0_144_1273 ();
 sg13g2_fill_8 FILLER_0_144_1281 ();
 sg13g2_fill_8 FILLER_0_144_1289 ();
 sg13g2_fill_8 FILLER_0_145_0 ();
 sg13g2_fill_8 FILLER_0_145_8 ();
 sg13g2_fill_8 FILLER_0_145_16 ();
 sg13g2_fill_8 FILLER_0_145_24 ();
 sg13g2_fill_8 FILLER_0_145_32 ();
 sg13g2_fill_8 FILLER_0_145_40 ();
 sg13g2_fill_8 FILLER_0_145_48 ();
 sg13g2_fill_8 FILLER_0_145_56 ();
 sg13g2_fill_8 FILLER_0_145_64 ();
 sg13g2_fill_8 FILLER_0_145_72 ();
 sg13g2_fill_8 FILLER_0_145_80 ();
 sg13g2_fill_8 FILLER_0_145_88 ();
 sg13g2_fill_8 FILLER_0_145_96 ();
 sg13g2_fill_8 FILLER_0_145_104 ();
 sg13g2_fill_8 FILLER_0_145_112 ();
 sg13g2_fill_8 FILLER_0_145_120 ();
 sg13g2_fill_8 FILLER_0_145_128 ();
 sg13g2_fill_8 FILLER_0_145_136 ();
 sg13g2_fill_8 FILLER_0_145_144 ();
 sg13g2_fill_8 FILLER_0_145_152 ();
 sg13g2_fill_8 FILLER_0_145_160 ();
 sg13g2_fill_8 FILLER_0_145_168 ();
 sg13g2_fill_8 FILLER_0_145_176 ();
 sg13g2_fill_8 FILLER_0_145_184 ();
 sg13g2_fill_8 FILLER_0_145_192 ();
 sg13g2_fill_8 FILLER_0_145_200 ();
 sg13g2_fill_8 FILLER_0_145_208 ();
 sg13g2_fill_8 FILLER_0_145_216 ();
 sg13g2_fill_8 FILLER_0_145_224 ();
 sg13g2_fill_8 FILLER_0_145_232 ();
 sg13g2_fill_8 FILLER_0_145_240 ();
 sg13g2_fill_8 FILLER_0_145_248 ();
 sg13g2_fill_8 FILLER_0_145_256 ();
 sg13g2_fill_8 FILLER_0_145_264 ();
 sg13g2_fill_2 FILLER_0_145_272 ();
 sg13g2_fill_1 FILLER_0_145_274 ();
 sg13g2_fill_2 FILLER_0_145_301 ();
 sg13g2_fill_4 FILLER_0_145_308 ();
 sg13g2_fill_4 FILLER_0_145_333 ();
 sg13g2_fill_2 FILLER_0_145_337 ();
 sg13g2_fill_4 FILLER_0_145_365 ();
 sg13g2_fill_2 FILLER_0_145_369 ();
 sg13g2_fill_4 FILLER_0_145_376 ();
 sg13g2_fill_2 FILLER_0_145_380 ();
 sg13g2_fill_8 FILLER_0_145_387 ();
 sg13g2_fill_2 FILLER_0_145_395 ();
 sg13g2_fill_1 FILLER_0_145_397 ();
 sg13g2_fill_2 FILLER_0_145_403 ();
 sg13g2_fill_2 FILLER_0_145_409 ();
 sg13g2_fill_8 FILLER_0_145_415 ();
 sg13g2_fill_8 FILLER_0_145_423 ();
 sg13g2_fill_8 FILLER_0_145_431 ();
 sg13g2_fill_2 FILLER_0_145_439 ();
 sg13g2_fill_1 FILLER_0_145_441 ();
 sg13g2_fill_8 FILLER_0_145_446 ();
 sg13g2_fill_8 FILLER_0_145_454 ();
 sg13g2_fill_8 FILLER_0_145_462 ();
 sg13g2_fill_8 FILLER_0_145_470 ();
 sg13g2_fill_8 FILLER_0_145_478 ();
 sg13g2_fill_8 FILLER_0_145_486 ();
 sg13g2_fill_8 FILLER_0_145_494 ();
 sg13g2_fill_8 FILLER_0_145_502 ();
 sg13g2_fill_8 FILLER_0_145_516 ();
 sg13g2_fill_2 FILLER_0_145_524 ();
 sg13g2_fill_2 FILLER_0_145_552 ();
 sg13g2_fill_8 FILLER_0_145_558 ();
 sg13g2_fill_2 FILLER_0_145_566 ();
 sg13g2_fill_8 FILLER_0_145_594 ();
 sg13g2_fill_4 FILLER_0_145_602 ();
 sg13g2_fill_2 FILLER_0_145_606 ();
 sg13g2_fill_1 FILLER_0_145_608 ();
 sg13g2_fill_2 FILLER_0_145_613 ();
 sg13g2_fill_2 FILLER_0_145_620 ();
 sg13g2_fill_2 FILLER_0_145_626 ();
 sg13g2_fill_8 FILLER_0_145_633 ();
 sg13g2_fill_8 FILLER_0_145_645 ();
 sg13g2_fill_8 FILLER_0_145_653 ();
 sg13g2_fill_4 FILLER_0_145_661 ();
 sg13g2_fill_1 FILLER_0_145_665 ();
 sg13g2_fill_2 FILLER_0_145_674 ();
 sg13g2_fill_4 FILLER_0_145_680 ();
 sg13g2_fill_2 FILLER_0_145_684 ();
 sg13g2_fill_1 FILLER_0_145_686 ();
 sg13g2_fill_8 FILLER_0_145_693 ();
 sg13g2_fill_8 FILLER_0_145_701 ();
 sg13g2_fill_8 FILLER_0_145_709 ();
 sg13g2_fill_8 FILLER_0_145_717 ();
 sg13g2_fill_1 FILLER_0_145_725 ();
 sg13g2_fill_2 FILLER_0_145_730 ();
 sg13g2_fill_4 FILLER_0_145_736 ();
 sg13g2_fill_2 FILLER_0_145_746 ();
 sg13g2_fill_2 FILLER_0_145_753 ();
 sg13g2_fill_2 FILLER_0_145_781 ();
 sg13g2_fill_8 FILLER_0_145_787 ();
 sg13g2_fill_8 FILLER_0_145_795 ();
 sg13g2_fill_4 FILLER_0_145_803 ();
 sg13g2_fill_2 FILLER_0_145_807 ();
 sg13g2_fill_4 FILLER_0_145_813 ();
 sg13g2_fill_2 FILLER_0_145_817 ();
 sg13g2_fill_2 FILLER_0_145_823 ();
 sg13g2_fill_8 FILLER_0_145_851 ();
 sg13g2_fill_8 FILLER_0_145_859 ();
 sg13g2_fill_8 FILLER_0_145_893 ();
 sg13g2_fill_8 FILLER_0_145_901 ();
 sg13g2_fill_2 FILLER_0_145_909 ();
 sg13g2_fill_2 FILLER_0_145_916 ();
 sg13g2_fill_8 FILLER_0_145_922 ();
 sg13g2_fill_8 FILLER_0_145_930 ();
 sg13g2_fill_4 FILLER_0_145_938 ();
 sg13g2_fill_2 FILLER_0_145_942 ();
 sg13g2_fill_1 FILLER_0_145_944 ();
 sg13g2_fill_8 FILLER_0_145_971 ();
 sg13g2_fill_8 FILLER_0_145_984 ();
 sg13g2_fill_8 FILLER_0_145_992 ();
 sg13g2_fill_4 FILLER_0_145_1000 ();
 sg13g2_fill_1 FILLER_0_145_1004 ();
 sg13g2_fill_2 FILLER_0_145_1012 ();
 sg13g2_fill_8 FILLER_0_145_1019 ();
 sg13g2_fill_8 FILLER_0_145_1027 ();
 sg13g2_fill_8 FILLER_0_145_1035 ();
 sg13g2_fill_8 FILLER_0_145_1043 ();
 sg13g2_fill_8 FILLER_0_145_1051 ();
 sg13g2_fill_2 FILLER_0_145_1059 ();
 sg13g2_fill_2 FILLER_0_145_1066 ();
 sg13g2_fill_2 FILLER_0_145_1094 ();
 sg13g2_fill_2 FILLER_0_145_1101 ();
 sg13g2_fill_1 FILLER_0_145_1103 ();
 sg13g2_fill_2 FILLER_0_145_1109 ();
 sg13g2_fill_1 FILLER_0_145_1111 ();
 sg13g2_fill_2 FILLER_0_145_1138 ();
 sg13g2_fill_8 FILLER_0_145_1145 ();
 sg13g2_fill_8 FILLER_0_145_1153 ();
 sg13g2_fill_8 FILLER_0_145_1161 ();
 sg13g2_fill_8 FILLER_0_145_1169 ();
 sg13g2_fill_2 FILLER_0_145_1177 ();
 sg13g2_fill_2 FILLER_0_145_1183 ();
 sg13g2_fill_2 FILLER_0_145_1190 ();
 sg13g2_fill_1 FILLER_0_145_1192 ();
 sg13g2_fill_2 FILLER_0_145_1219 ();
 sg13g2_fill_1 FILLER_0_145_1221 ();
 sg13g2_fill_4 FILLER_0_145_1226 ();
 sg13g2_fill_2 FILLER_0_145_1235 ();
 sg13g2_fill_4 FILLER_0_145_1242 ();
 sg13g2_fill_2 FILLER_0_145_1246 ();
 sg13g2_fill_1 FILLER_0_145_1248 ();
 sg13g2_fill_8 FILLER_0_145_1253 ();
 sg13g2_fill_8 FILLER_0_145_1261 ();
 sg13g2_fill_8 FILLER_0_145_1269 ();
 sg13g2_fill_8 FILLER_0_145_1277 ();
 sg13g2_fill_8 FILLER_0_145_1285 ();
 sg13g2_fill_4 FILLER_0_145_1293 ();
 sg13g2_fill_8 FILLER_0_146_0 ();
 sg13g2_fill_8 FILLER_0_146_8 ();
 sg13g2_fill_8 FILLER_0_146_16 ();
 sg13g2_fill_8 FILLER_0_146_24 ();
 sg13g2_fill_8 FILLER_0_146_32 ();
 sg13g2_fill_8 FILLER_0_146_40 ();
 sg13g2_fill_8 FILLER_0_146_48 ();
 sg13g2_fill_8 FILLER_0_146_56 ();
 sg13g2_fill_8 FILLER_0_146_64 ();
 sg13g2_fill_8 FILLER_0_146_72 ();
 sg13g2_fill_8 FILLER_0_146_80 ();
 sg13g2_fill_8 FILLER_0_146_88 ();
 sg13g2_fill_8 FILLER_0_146_96 ();
 sg13g2_fill_8 FILLER_0_146_104 ();
 sg13g2_fill_8 FILLER_0_146_112 ();
 sg13g2_fill_8 FILLER_0_146_120 ();
 sg13g2_fill_8 FILLER_0_146_128 ();
 sg13g2_fill_8 FILLER_0_146_136 ();
 sg13g2_fill_8 FILLER_0_146_144 ();
 sg13g2_fill_8 FILLER_0_146_152 ();
 sg13g2_fill_8 FILLER_0_146_160 ();
 sg13g2_fill_8 FILLER_0_146_168 ();
 sg13g2_fill_8 FILLER_0_146_176 ();
 sg13g2_fill_8 FILLER_0_146_184 ();
 sg13g2_fill_8 FILLER_0_146_192 ();
 sg13g2_fill_8 FILLER_0_146_200 ();
 sg13g2_fill_8 FILLER_0_146_208 ();
 sg13g2_fill_8 FILLER_0_146_216 ();
 sg13g2_fill_8 FILLER_0_146_224 ();
 sg13g2_fill_8 FILLER_0_146_232 ();
 sg13g2_fill_8 FILLER_0_146_240 ();
 sg13g2_fill_8 FILLER_0_146_248 ();
 sg13g2_fill_8 FILLER_0_146_256 ();
 sg13g2_fill_8 FILLER_0_146_264 ();
 sg13g2_fill_2 FILLER_0_146_272 ();
 sg13g2_fill_1 FILLER_0_146_274 ();
 sg13g2_fill_2 FILLER_0_146_301 ();
 sg13g2_fill_8 FILLER_0_146_329 ();
 sg13g2_fill_4 FILLER_0_146_337 ();
 sg13g2_fill_2 FILLER_0_146_341 ();
 sg13g2_fill_4 FILLER_0_146_348 ();
 sg13g2_fill_2 FILLER_0_146_378 ();
 sg13g2_fill_8 FILLER_0_146_385 ();
 sg13g2_fill_8 FILLER_0_146_419 ();
 sg13g2_fill_8 FILLER_0_146_427 ();
 sg13g2_fill_8 FILLER_0_146_435 ();
 sg13g2_fill_4 FILLER_0_146_443 ();
 sg13g2_fill_8 FILLER_0_146_452 ();
 sg13g2_fill_8 FILLER_0_146_460 ();
 sg13g2_fill_8 FILLER_0_146_468 ();
 sg13g2_fill_1 FILLER_0_146_476 ();
 sg13g2_fill_8 FILLER_0_146_482 ();
 sg13g2_fill_8 FILLER_0_146_490 ();
 sg13g2_fill_1 FILLER_0_146_498 ();
 sg13g2_fill_8 FILLER_0_146_509 ();
 sg13g2_fill_8 FILLER_0_146_517 ();
 sg13g2_fill_4 FILLER_0_146_525 ();
 sg13g2_fill_2 FILLER_0_146_529 ();
 sg13g2_fill_8 FILLER_0_146_536 ();
 sg13g2_fill_8 FILLER_0_146_544 ();
 sg13g2_fill_8 FILLER_0_146_552 ();
 sg13g2_fill_2 FILLER_0_146_560 ();
 sg13g2_fill_8 FILLER_0_146_583 ();
 sg13g2_fill_8 FILLER_0_146_591 ();
 sg13g2_fill_4 FILLER_0_146_599 ();
 sg13g2_fill_2 FILLER_0_146_603 ();
 sg13g2_fill_1 FILLER_0_146_605 ();
 sg13g2_fill_8 FILLER_0_146_611 ();
 sg13g2_fill_8 FILLER_0_146_619 ();
 sg13g2_fill_8 FILLER_0_146_627 ();
 sg13g2_fill_8 FILLER_0_146_635 ();
 sg13g2_fill_8 FILLER_0_146_643 ();
 sg13g2_fill_8 FILLER_0_146_651 ();
 sg13g2_fill_8 FILLER_0_146_659 ();
 sg13g2_fill_2 FILLER_0_146_667 ();
 sg13g2_fill_1 FILLER_0_146_669 ();
 sg13g2_fill_8 FILLER_0_146_675 ();
 sg13g2_fill_8 FILLER_0_146_683 ();
 sg13g2_fill_8 FILLER_0_146_691 ();
 sg13g2_fill_4 FILLER_0_146_699 ();
 sg13g2_fill_8 FILLER_0_146_708 ();
 sg13g2_fill_4 FILLER_0_146_716 ();
 sg13g2_fill_2 FILLER_0_146_720 ();
 sg13g2_fill_1 FILLER_0_146_722 ();
 sg13g2_fill_4 FILLER_0_146_729 ();
 sg13g2_fill_1 FILLER_0_146_733 ();
 sg13g2_fill_4 FILLER_0_146_740 ();
 sg13g2_fill_2 FILLER_0_146_748 ();
 sg13g2_fill_4 FILLER_0_146_758 ();
 sg13g2_fill_2 FILLER_0_146_762 ();
 sg13g2_fill_2 FILLER_0_146_769 ();
 sg13g2_fill_8 FILLER_0_146_776 ();
 sg13g2_fill_8 FILLER_0_146_784 ();
 sg13g2_fill_8 FILLER_0_146_792 ();
 sg13g2_fill_8 FILLER_0_146_800 ();
 sg13g2_fill_1 FILLER_0_146_808 ();
 sg13g2_fill_2 FILLER_0_146_814 ();
 sg13g2_fill_2 FILLER_0_146_842 ();
 sg13g2_fill_2 FILLER_0_146_849 ();
 sg13g2_fill_8 FILLER_0_146_857 ();
 sg13g2_fill_8 FILLER_0_146_865 ();
 sg13g2_fill_8 FILLER_0_146_873 ();
 sg13g2_fill_8 FILLER_0_146_881 ();
 sg13g2_fill_8 FILLER_0_146_889 ();
 sg13g2_fill_8 FILLER_0_146_897 ();
 sg13g2_fill_8 FILLER_0_146_905 ();
 sg13g2_fill_8 FILLER_0_146_913 ();
 sg13g2_fill_8 FILLER_0_146_921 ();
 sg13g2_fill_4 FILLER_0_146_929 ();
 sg13g2_fill_2 FILLER_0_146_933 ();
 sg13g2_fill_2 FILLER_0_146_940 ();
 sg13g2_fill_2 FILLER_0_146_946 ();
 sg13g2_fill_1 FILLER_0_146_948 ();
 sg13g2_fill_4 FILLER_0_146_970 ();
 sg13g2_fill_4 FILLER_0_146_978 ();
 sg13g2_fill_4 FILLER_0_146_1008 ();
 sg13g2_fill_1 FILLER_0_146_1012 ();
 sg13g2_fill_8 FILLER_0_146_1017 ();
 sg13g2_fill_4 FILLER_0_146_1025 ();
 sg13g2_fill_1 FILLER_0_146_1029 ();
 sg13g2_fill_2 FILLER_0_146_1035 ();
 sg13g2_fill_2 FILLER_0_146_1041 ();
 sg13g2_fill_1 FILLER_0_146_1043 ();
 sg13g2_fill_8 FILLER_0_146_1054 ();
 sg13g2_fill_8 FILLER_0_146_1062 ();
 sg13g2_fill_8 FILLER_0_146_1070 ();
 sg13g2_fill_4 FILLER_0_146_1083 ();
 sg13g2_fill_4 FILLER_0_146_1091 ();
 sg13g2_fill_1 FILLER_0_146_1095 ();
 sg13g2_fill_4 FILLER_0_146_1102 ();
 sg13g2_fill_4 FILLER_0_146_1114 ();
 sg13g2_fill_4 FILLER_0_146_1122 ();
 sg13g2_fill_1 FILLER_0_146_1126 ();
 sg13g2_fill_4 FILLER_0_146_1132 ();
 sg13g2_fill_2 FILLER_0_146_1136 ();
 sg13g2_fill_8 FILLER_0_146_1146 ();
 sg13g2_fill_8 FILLER_0_146_1154 ();
 sg13g2_fill_8 FILLER_0_146_1162 ();
 sg13g2_fill_8 FILLER_0_146_1170 ();
 sg13g2_fill_8 FILLER_0_146_1178 ();
 sg13g2_fill_8 FILLER_0_146_1186 ();
 sg13g2_fill_8 FILLER_0_146_1194 ();
 sg13g2_fill_8 FILLER_0_146_1202 ();
 sg13g2_fill_8 FILLER_0_146_1210 ();
 sg13g2_fill_8 FILLER_0_146_1218 ();
 sg13g2_fill_8 FILLER_0_146_1226 ();
 sg13g2_fill_8 FILLER_0_146_1234 ();
 sg13g2_fill_8 FILLER_0_146_1242 ();
 sg13g2_fill_8 FILLER_0_146_1250 ();
 sg13g2_fill_8 FILLER_0_146_1258 ();
 sg13g2_fill_8 FILLER_0_146_1266 ();
 sg13g2_fill_8 FILLER_0_146_1274 ();
 sg13g2_fill_8 FILLER_0_146_1282 ();
 sg13g2_fill_4 FILLER_0_146_1290 ();
 sg13g2_fill_2 FILLER_0_146_1294 ();
 sg13g2_fill_1 FILLER_0_146_1296 ();
 sg13g2_fill_8 FILLER_0_147_0 ();
 sg13g2_fill_8 FILLER_0_147_8 ();
 sg13g2_fill_8 FILLER_0_147_16 ();
 sg13g2_fill_8 FILLER_0_147_24 ();
 sg13g2_fill_8 FILLER_0_147_32 ();
 sg13g2_fill_8 FILLER_0_147_40 ();
 sg13g2_fill_8 FILLER_0_147_48 ();
 sg13g2_fill_8 FILLER_0_147_56 ();
 sg13g2_fill_8 FILLER_0_147_64 ();
 sg13g2_fill_8 FILLER_0_147_72 ();
 sg13g2_fill_8 FILLER_0_147_80 ();
 sg13g2_fill_8 FILLER_0_147_88 ();
 sg13g2_fill_8 FILLER_0_147_96 ();
 sg13g2_fill_8 FILLER_0_147_104 ();
 sg13g2_fill_8 FILLER_0_147_112 ();
 sg13g2_fill_8 FILLER_0_147_120 ();
 sg13g2_fill_8 FILLER_0_147_128 ();
 sg13g2_fill_8 FILLER_0_147_136 ();
 sg13g2_fill_8 FILLER_0_147_144 ();
 sg13g2_fill_8 FILLER_0_147_152 ();
 sg13g2_fill_8 FILLER_0_147_160 ();
 sg13g2_fill_8 FILLER_0_147_168 ();
 sg13g2_fill_8 FILLER_0_147_176 ();
 sg13g2_fill_8 FILLER_0_147_184 ();
 sg13g2_fill_8 FILLER_0_147_192 ();
 sg13g2_fill_8 FILLER_0_147_200 ();
 sg13g2_fill_8 FILLER_0_147_208 ();
 sg13g2_fill_8 FILLER_0_147_216 ();
 sg13g2_fill_8 FILLER_0_147_224 ();
 sg13g2_fill_8 FILLER_0_147_232 ();
 sg13g2_fill_8 FILLER_0_147_240 ();
 sg13g2_fill_8 FILLER_0_147_248 ();
 sg13g2_fill_8 FILLER_0_147_256 ();
 sg13g2_fill_8 FILLER_0_147_264 ();
 sg13g2_fill_2 FILLER_0_147_277 ();
 sg13g2_fill_2 FILLER_0_147_284 ();
 sg13g2_fill_2 FILLER_0_147_290 ();
 sg13g2_fill_1 FILLER_0_147_292 ();
 sg13g2_fill_4 FILLER_0_147_297 ();
 sg13g2_fill_2 FILLER_0_147_305 ();
 sg13g2_fill_8 FILLER_0_147_328 ();
 sg13g2_fill_1 FILLER_0_147_336 ();
 sg13g2_fill_2 FILLER_0_147_342 ();
 sg13g2_fill_4 FILLER_0_147_348 ();
 sg13g2_fill_4 FILLER_0_147_357 ();
 sg13g2_fill_1 FILLER_0_147_361 ();
 sg13g2_fill_2 FILLER_0_147_367 ();
 sg13g2_fill_2 FILLER_0_147_374 ();
 sg13g2_fill_2 FILLER_0_147_383 ();
 sg13g2_fill_1 FILLER_0_147_385 ();
 sg13g2_fill_2 FILLER_0_147_391 ();
 sg13g2_fill_4 FILLER_0_147_399 ();
 sg13g2_fill_1 FILLER_0_147_403 ();
 sg13g2_fill_8 FILLER_0_147_408 ();
 sg13g2_fill_8 FILLER_0_147_416 ();
 sg13g2_fill_8 FILLER_0_147_424 ();
 sg13g2_fill_8 FILLER_0_147_432 ();
 sg13g2_fill_8 FILLER_0_147_440 ();
 sg13g2_fill_8 FILLER_0_147_448 ();
 sg13g2_fill_8 FILLER_0_147_456 ();
 sg13g2_fill_8 FILLER_0_147_464 ();
 sg13g2_fill_2 FILLER_0_147_472 ();
 sg13g2_fill_2 FILLER_0_147_479 ();
 sg13g2_fill_1 FILLER_0_147_481 ();
 sg13g2_fill_8 FILLER_0_147_486 ();
 sg13g2_fill_8 FILLER_0_147_494 ();
 sg13g2_fill_8 FILLER_0_147_502 ();
 sg13g2_fill_8 FILLER_0_147_510 ();
 sg13g2_fill_4 FILLER_0_147_518 ();
 sg13g2_fill_4 FILLER_0_147_527 ();
 sg13g2_fill_1 FILLER_0_147_531 ();
 sg13g2_fill_8 FILLER_0_147_558 ();
 sg13g2_fill_8 FILLER_0_147_566 ();
 sg13g2_fill_8 FILLER_0_147_574 ();
 sg13g2_fill_8 FILLER_0_147_582 ();
 sg13g2_fill_8 FILLER_0_147_590 ();
 sg13g2_fill_8 FILLER_0_147_598 ();
 sg13g2_fill_8 FILLER_0_147_606 ();
 sg13g2_fill_2 FILLER_0_147_614 ();
 sg13g2_fill_1 FILLER_0_147_616 ();
 sg13g2_fill_2 FILLER_0_147_622 ();
 sg13g2_fill_2 FILLER_0_147_629 ();
 sg13g2_fill_2 FILLER_0_147_636 ();
 sg13g2_fill_1 FILLER_0_147_638 ();
 sg13g2_fill_8 FILLER_0_147_644 ();
 sg13g2_fill_2 FILLER_0_147_657 ();
 sg13g2_fill_4 FILLER_0_147_663 ();
 sg13g2_fill_2 FILLER_0_147_667 ();
 sg13g2_fill_1 FILLER_0_147_669 ();
 sg13g2_fill_4 FILLER_0_147_674 ();
 sg13g2_fill_2 FILLER_0_147_678 ();
 sg13g2_fill_8 FILLER_0_147_685 ();
 sg13g2_fill_8 FILLER_0_147_693 ();
 sg13g2_fill_4 FILLER_0_147_701 ();
 sg13g2_fill_2 FILLER_0_147_705 ();
 sg13g2_fill_8 FILLER_0_147_712 ();
 sg13g2_fill_8 FILLER_0_147_720 ();
 sg13g2_fill_8 FILLER_0_147_728 ();
 sg13g2_fill_4 FILLER_0_147_736 ();
 sg13g2_fill_2 FILLER_0_147_740 ();
 sg13g2_fill_4 FILLER_0_147_747 ();
 sg13g2_fill_8 FILLER_0_147_756 ();
 sg13g2_fill_4 FILLER_0_147_764 ();
 sg13g2_fill_2 FILLER_0_147_768 ();
 sg13g2_fill_4 FILLER_0_147_778 ();
 sg13g2_fill_2 FILLER_0_147_782 ();
 sg13g2_fill_1 FILLER_0_147_784 ();
 sg13g2_fill_2 FILLER_0_147_790 ();
 sg13g2_fill_8 FILLER_0_147_802 ();
 sg13g2_fill_8 FILLER_0_147_810 ();
 sg13g2_fill_8 FILLER_0_147_818 ();
 sg13g2_fill_8 FILLER_0_147_826 ();
 sg13g2_fill_8 FILLER_0_147_834 ();
 sg13g2_fill_8 FILLER_0_147_842 ();
 sg13g2_fill_8 FILLER_0_147_850 ();
 sg13g2_fill_8 FILLER_0_147_858 ();
 sg13g2_fill_8 FILLER_0_147_866 ();
 sg13g2_fill_8 FILLER_0_147_874 ();
 sg13g2_fill_4 FILLER_0_147_882 ();
 sg13g2_fill_1 FILLER_0_147_886 ();
 sg13g2_fill_8 FILLER_0_147_892 ();
 sg13g2_fill_8 FILLER_0_147_900 ();
 sg13g2_fill_8 FILLER_0_147_908 ();
 sg13g2_fill_2 FILLER_0_147_919 ();
 sg13g2_fill_8 FILLER_0_147_947 ();
 sg13g2_fill_8 FILLER_0_147_955 ();
 sg13g2_fill_8 FILLER_0_147_963 ();
 sg13g2_fill_4 FILLER_0_147_971 ();
 sg13g2_fill_1 FILLER_0_147_975 ();
 sg13g2_fill_8 FILLER_0_147_983 ();
 sg13g2_fill_8 FILLER_0_147_991 ();
 sg13g2_fill_8 FILLER_0_147_999 ();
 sg13g2_fill_8 FILLER_0_147_1007 ();
 sg13g2_fill_8 FILLER_0_147_1015 ();
 sg13g2_fill_2 FILLER_0_147_1027 ();
 sg13g2_fill_4 FILLER_0_147_1055 ();
 sg13g2_fill_2 FILLER_0_147_1059 ();
 sg13g2_fill_8 FILLER_0_147_1066 ();
 sg13g2_fill_8 FILLER_0_147_1074 ();
 sg13g2_fill_8 FILLER_0_147_1082 ();
 sg13g2_fill_4 FILLER_0_147_1090 ();
 sg13g2_fill_1 FILLER_0_147_1094 ();
 sg13g2_fill_8 FILLER_0_147_1100 ();
 sg13g2_fill_1 FILLER_0_147_1108 ();
 sg13g2_fill_4 FILLER_0_147_1114 ();
 sg13g2_fill_2 FILLER_0_147_1118 ();
 sg13g2_fill_1 FILLER_0_147_1120 ();
 sg13g2_fill_8 FILLER_0_147_1125 ();
 sg13g2_fill_4 FILLER_0_147_1139 ();
 sg13g2_fill_8 FILLER_0_147_1148 ();
 sg13g2_fill_8 FILLER_0_147_1156 ();
 sg13g2_fill_8 FILLER_0_147_1164 ();
 sg13g2_fill_2 FILLER_0_147_1172 ();
 sg13g2_fill_8 FILLER_0_147_1184 ();
 sg13g2_fill_8 FILLER_0_147_1192 ();
 sg13g2_fill_8 FILLER_0_147_1200 ();
 sg13g2_fill_4 FILLER_0_147_1208 ();
 sg13g2_fill_4 FILLER_0_147_1233 ();
 sg13g2_fill_2 FILLER_0_147_1237 ();
 sg13g2_fill_8 FILLER_0_147_1249 ();
 sg13g2_fill_8 FILLER_0_147_1257 ();
 sg13g2_fill_8 FILLER_0_147_1265 ();
 sg13g2_fill_8 FILLER_0_147_1273 ();
 sg13g2_fill_8 FILLER_0_147_1281 ();
 sg13g2_fill_8 FILLER_0_147_1289 ();
 sg13g2_fill_8 FILLER_0_148_0 ();
 sg13g2_fill_8 FILLER_0_148_8 ();
 sg13g2_fill_8 FILLER_0_148_16 ();
 sg13g2_fill_8 FILLER_0_148_24 ();
 sg13g2_fill_8 FILLER_0_148_32 ();
 sg13g2_fill_8 FILLER_0_148_40 ();
 sg13g2_fill_8 FILLER_0_148_48 ();
 sg13g2_fill_8 FILLER_0_148_56 ();
 sg13g2_fill_8 FILLER_0_148_64 ();
 sg13g2_fill_8 FILLER_0_148_72 ();
 sg13g2_fill_8 FILLER_0_148_80 ();
 sg13g2_fill_8 FILLER_0_148_88 ();
 sg13g2_fill_8 FILLER_0_148_96 ();
 sg13g2_fill_8 FILLER_0_148_104 ();
 sg13g2_fill_8 FILLER_0_148_112 ();
 sg13g2_fill_8 FILLER_0_148_120 ();
 sg13g2_fill_8 FILLER_0_148_128 ();
 sg13g2_fill_8 FILLER_0_148_136 ();
 sg13g2_fill_8 FILLER_0_148_144 ();
 sg13g2_fill_8 FILLER_0_148_152 ();
 sg13g2_fill_8 FILLER_0_148_160 ();
 sg13g2_fill_8 FILLER_0_148_168 ();
 sg13g2_fill_8 FILLER_0_148_176 ();
 sg13g2_fill_8 FILLER_0_148_184 ();
 sg13g2_fill_8 FILLER_0_148_192 ();
 sg13g2_fill_8 FILLER_0_148_200 ();
 sg13g2_fill_8 FILLER_0_148_208 ();
 sg13g2_fill_8 FILLER_0_148_216 ();
 sg13g2_fill_8 FILLER_0_148_224 ();
 sg13g2_fill_8 FILLER_0_148_232 ();
 sg13g2_fill_8 FILLER_0_148_240 ();
 sg13g2_fill_8 FILLER_0_148_248 ();
 sg13g2_fill_8 FILLER_0_148_256 ();
 sg13g2_fill_8 FILLER_0_148_264 ();
 sg13g2_fill_8 FILLER_0_148_272 ();
 sg13g2_fill_8 FILLER_0_148_280 ();
 sg13g2_fill_8 FILLER_0_148_288 ();
 sg13g2_fill_8 FILLER_0_148_296 ();
 sg13g2_fill_8 FILLER_0_148_304 ();
 sg13g2_fill_8 FILLER_0_148_312 ();
 sg13g2_fill_8 FILLER_0_148_320 ();
 sg13g2_fill_8 FILLER_0_148_328 ();
 sg13g2_fill_8 FILLER_0_148_336 ();
 sg13g2_fill_4 FILLER_0_148_344 ();
 sg13g2_fill_1 FILLER_0_148_348 ();
 sg13g2_fill_8 FILLER_0_148_370 ();
 sg13g2_fill_4 FILLER_0_148_378 ();
 sg13g2_fill_2 FILLER_0_148_382 ();
 sg13g2_fill_1 FILLER_0_148_384 ();
 sg13g2_fill_8 FILLER_0_148_389 ();
 sg13g2_fill_8 FILLER_0_148_397 ();
 sg13g2_fill_8 FILLER_0_148_405 ();
 sg13g2_fill_8 FILLER_0_148_413 ();
 sg13g2_fill_4 FILLER_0_148_421 ();
 sg13g2_fill_2 FILLER_0_148_425 ();
 sg13g2_fill_1 FILLER_0_148_427 ();
 sg13g2_fill_8 FILLER_0_148_433 ();
 sg13g2_fill_8 FILLER_0_148_441 ();
 sg13g2_fill_8 FILLER_0_148_449 ();
 sg13g2_fill_4 FILLER_0_148_457 ();
 sg13g2_fill_8 FILLER_0_148_466 ();
 sg13g2_fill_2 FILLER_0_148_474 ();
 sg13g2_fill_4 FILLER_0_148_502 ();
 sg13g2_fill_1 FILLER_0_148_506 ();
 sg13g2_fill_8 FILLER_0_148_512 ();
 sg13g2_fill_8 FILLER_0_148_520 ();
 sg13g2_fill_2 FILLER_0_148_528 ();
 sg13g2_fill_1 FILLER_0_148_530 ();
 sg13g2_fill_8 FILLER_0_148_536 ();
 sg13g2_fill_8 FILLER_0_148_544 ();
 sg13g2_fill_1 FILLER_0_148_552 ();
 sg13g2_fill_8 FILLER_0_148_574 ();
 sg13g2_fill_8 FILLER_0_148_582 ();
 sg13g2_fill_8 FILLER_0_148_590 ();
 sg13g2_fill_8 FILLER_0_148_598 ();
 sg13g2_fill_8 FILLER_0_148_606 ();
 sg13g2_fill_8 FILLER_0_148_614 ();
 sg13g2_fill_1 FILLER_0_148_622 ();
 sg13g2_fill_8 FILLER_0_148_628 ();
 sg13g2_fill_4 FILLER_0_148_636 ();
 sg13g2_fill_2 FILLER_0_148_646 ();
 sg13g2_fill_2 FILLER_0_148_674 ();
 sg13g2_fill_2 FILLER_0_148_680 ();
 sg13g2_fill_4 FILLER_0_148_708 ();
 sg13g2_fill_8 FILLER_0_148_717 ();
 sg13g2_fill_8 FILLER_0_148_725 ();
 sg13g2_fill_4 FILLER_0_148_733 ();
 sg13g2_fill_2 FILLER_0_148_737 ();
 sg13g2_fill_8 FILLER_0_148_765 ();
 sg13g2_fill_1 FILLER_0_148_773 ();
 sg13g2_fill_2 FILLER_0_148_779 ();
 sg13g2_fill_8 FILLER_0_148_807 ();
 sg13g2_fill_8 FILLER_0_148_815 ();
 sg13g2_fill_4 FILLER_0_148_823 ();
 sg13g2_fill_2 FILLER_0_148_827 ();
 sg13g2_fill_1 FILLER_0_148_829 ();
 sg13g2_fill_2 FILLER_0_148_835 ();
 sg13g2_fill_8 FILLER_0_148_842 ();
 sg13g2_fill_1 FILLER_0_148_850 ();
 sg13g2_fill_4 FILLER_0_148_855 ();
 sg13g2_fill_2 FILLER_0_148_864 ();
 sg13g2_fill_2 FILLER_0_148_870 ();
 sg13g2_fill_2 FILLER_0_148_893 ();
 sg13g2_fill_4 FILLER_0_148_899 ();
 sg13g2_fill_2 FILLER_0_148_903 ();
 sg13g2_fill_2 FILLER_0_148_910 ();
 sg13g2_fill_8 FILLER_0_148_918 ();
 sg13g2_fill_8 FILLER_0_148_926 ();
 sg13g2_fill_8 FILLER_0_148_934 ();
 sg13g2_fill_4 FILLER_0_148_942 ();
 sg13g2_fill_2 FILLER_0_148_946 ();
 sg13g2_fill_1 FILLER_0_148_948 ();
 sg13g2_fill_8 FILLER_0_148_954 ();
 sg13g2_fill_8 FILLER_0_148_962 ();
 sg13g2_fill_8 FILLER_0_148_970 ();
 sg13g2_fill_4 FILLER_0_148_978 ();
 sg13g2_fill_1 FILLER_0_148_982 ();
 sg13g2_fill_4 FILLER_0_148_989 ();
 sg13g2_fill_2 FILLER_0_148_993 ();
 sg13g2_fill_2 FILLER_0_148_1021 ();
 sg13g2_fill_8 FILLER_0_148_1028 ();
 sg13g2_fill_8 FILLER_0_148_1036 ();
 sg13g2_fill_8 FILLER_0_148_1044 ();
 sg13g2_fill_4 FILLER_0_148_1052 ();
 sg13g2_fill_8 FILLER_0_148_1061 ();
 sg13g2_fill_4 FILLER_0_148_1069 ();
 sg13g2_fill_2 FILLER_0_148_1073 ();
 sg13g2_fill_1 FILLER_0_148_1075 ();
 sg13g2_fill_8 FILLER_0_148_1081 ();
 sg13g2_fill_8 FILLER_0_148_1089 ();
 sg13g2_fill_8 FILLER_0_148_1097 ();
 sg13g2_fill_2 FILLER_0_148_1105 ();
 sg13g2_fill_8 FILLER_0_148_1112 ();
 sg13g2_fill_8 FILLER_0_148_1120 ();
 sg13g2_fill_8 FILLER_0_148_1128 ();
 sg13g2_fill_8 FILLER_0_148_1136 ();
 sg13g2_fill_8 FILLER_0_148_1144 ();
 sg13g2_fill_8 FILLER_0_148_1152 ();
 sg13g2_fill_8 FILLER_0_148_1160 ();
 sg13g2_fill_2 FILLER_0_148_1168 ();
 sg13g2_fill_2 FILLER_0_148_1174 ();
 sg13g2_fill_4 FILLER_0_148_1180 ();
 sg13g2_fill_2 FILLER_0_148_1188 ();
 sg13g2_fill_2 FILLER_0_148_1216 ();
 sg13g2_fill_8 FILLER_0_148_1244 ();
 sg13g2_fill_8 FILLER_0_148_1252 ();
 sg13g2_fill_8 FILLER_0_148_1260 ();
 sg13g2_fill_8 FILLER_0_148_1268 ();
 sg13g2_fill_8 FILLER_0_148_1276 ();
 sg13g2_fill_8 FILLER_0_148_1284 ();
 sg13g2_fill_4 FILLER_0_148_1292 ();
 sg13g2_fill_1 FILLER_0_148_1296 ();
 sg13g2_fill_8 FILLER_0_149_0 ();
 sg13g2_fill_8 FILLER_0_149_8 ();
 sg13g2_fill_8 FILLER_0_149_16 ();
 sg13g2_fill_8 FILLER_0_149_24 ();
 sg13g2_fill_8 FILLER_0_149_32 ();
 sg13g2_fill_8 FILLER_0_149_40 ();
 sg13g2_fill_8 FILLER_0_149_48 ();
 sg13g2_fill_8 FILLER_0_149_56 ();
 sg13g2_fill_8 FILLER_0_149_64 ();
 sg13g2_fill_8 FILLER_0_149_72 ();
 sg13g2_fill_8 FILLER_0_149_80 ();
 sg13g2_fill_8 FILLER_0_149_88 ();
 sg13g2_fill_8 FILLER_0_149_96 ();
 sg13g2_fill_8 FILLER_0_149_104 ();
 sg13g2_fill_8 FILLER_0_149_112 ();
 sg13g2_fill_8 FILLER_0_149_120 ();
 sg13g2_fill_8 FILLER_0_149_128 ();
 sg13g2_fill_8 FILLER_0_149_136 ();
 sg13g2_fill_8 FILLER_0_149_144 ();
 sg13g2_fill_8 FILLER_0_149_152 ();
 sg13g2_fill_8 FILLER_0_149_160 ();
 sg13g2_fill_8 FILLER_0_149_168 ();
 sg13g2_fill_8 FILLER_0_149_176 ();
 sg13g2_fill_8 FILLER_0_149_184 ();
 sg13g2_fill_8 FILLER_0_149_192 ();
 sg13g2_fill_8 FILLER_0_149_200 ();
 sg13g2_fill_8 FILLER_0_149_208 ();
 sg13g2_fill_8 FILLER_0_149_216 ();
 sg13g2_fill_8 FILLER_0_149_224 ();
 sg13g2_fill_8 FILLER_0_149_232 ();
 sg13g2_fill_8 FILLER_0_149_240 ();
 sg13g2_fill_8 FILLER_0_149_248 ();
 sg13g2_fill_8 FILLER_0_149_256 ();
 sg13g2_fill_8 FILLER_0_149_264 ();
 sg13g2_fill_8 FILLER_0_149_272 ();
 sg13g2_fill_8 FILLER_0_149_280 ();
 sg13g2_fill_8 FILLER_0_149_288 ();
 sg13g2_fill_8 FILLER_0_149_296 ();
 sg13g2_fill_8 FILLER_0_149_304 ();
 sg13g2_fill_8 FILLER_0_149_312 ();
 sg13g2_fill_2 FILLER_0_149_320 ();
 sg13g2_fill_1 FILLER_0_149_322 ();
 sg13g2_fill_8 FILLER_0_149_328 ();
 sg13g2_fill_1 FILLER_0_149_336 ();
 sg13g2_fill_8 FILLER_0_149_342 ();
 sg13g2_fill_8 FILLER_0_149_350 ();
 sg13g2_fill_8 FILLER_0_149_358 ();
 sg13g2_fill_4 FILLER_0_149_366 ();
 sg13g2_fill_2 FILLER_0_149_370 ();
 sg13g2_fill_8 FILLER_0_149_375 ();
 sg13g2_fill_4 FILLER_0_149_383 ();
 sg13g2_fill_8 FILLER_0_149_392 ();
 sg13g2_fill_2 FILLER_0_149_400 ();
 sg13g2_fill_8 FILLER_0_149_407 ();
 sg13g2_fill_1 FILLER_0_149_415 ();
 sg13g2_fill_2 FILLER_0_149_421 ();
 sg13g2_fill_8 FILLER_0_149_427 ();
 sg13g2_fill_4 FILLER_0_149_435 ();
 sg13g2_fill_2 FILLER_0_149_439 ();
 sg13g2_fill_2 FILLER_0_149_467 ();
 sg13g2_fill_4 FILLER_0_149_473 ();
 sg13g2_fill_2 FILLER_0_149_477 ();
 sg13g2_fill_1 FILLER_0_149_479 ();
 sg13g2_fill_8 FILLER_0_149_501 ();
 sg13g2_fill_8 FILLER_0_149_509 ();
 sg13g2_fill_2 FILLER_0_149_517 ();
 sg13g2_fill_1 FILLER_0_149_519 ();
 sg13g2_fill_8 FILLER_0_149_525 ();
 sg13g2_fill_4 FILLER_0_149_533 ();
 sg13g2_fill_2 FILLER_0_149_541 ();
 sg13g2_fill_2 FILLER_0_149_548 ();
 sg13g2_fill_8 FILLER_0_149_555 ();
 sg13g2_fill_8 FILLER_0_149_563 ();
 sg13g2_fill_1 FILLER_0_149_571 ();
 sg13g2_fill_2 FILLER_0_149_576 ();
 sg13g2_fill_2 FILLER_0_149_583 ();
 sg13g2_fill_2 FILLER_0_149_589 ();
 sg13g2_fill_2 FILLER_0_149_617 ();
 sg13g2_fill_1 FILLER_0_149_619 ();
 sg13g2_fill_2 FILLER_0_149_646 ();
 sg13g2_fill_1 FILLER_0_149_648 ();
 sg13g2_fill_4 FILLER_0_149_654 ();
 sg13g2_fill_4 FILLER_0_149_666 ();
 sg13g2_fill_4 FILLER_0_149_676 ();
 sg13g2_fill_1 FILLER_0_149_680 ();
 sg13g2_fill_2 FILLER_0_149_686 ();
 sg13g2_fill_2 FILLER_0_149_709 ();
 sg13g2_fill_8 FILLER_0_149_715 ();
 sg13g2_fill_8 FILLER_0_149_723 ();
 sg13g2_fill_8 FILLER_0_149_731 ();
 sg13g2_fill_8 FILLER_0_149_739 ();
 sg13g2_fill_8 FILLER_0_149_747 ();
 sg13g2_fill_4 FILLER_0_149_755 ();
 sg13g2_fill_2 FILLER_0_149_759 ();
 sg13g2_fill_2 FILLER_0_149_766 ();
 sg13g2_fill_4 FILLER_0_149_773 ();
 sg13g2_fill_2 FILLER_0_149_777 ();
 sg13g2_fill_1 FILLER_0_149_779 ();
 sg13g2_fill_8 FILLER_0_149_784 ();
 sg13g2_fill_8 FILLER_0_149_818 ();
 sg13g2_fill_2 FILLER_0_149_826 ();
 sg13g2_fill_1 FILLER_0_149_828 ();
 sg13g2_fill_4 FILLER_0_149_834 ();
 sg13g2_fill_2 FILLER_0_149_838 ();
 sg13g2_fill_1 FILLER_0_149_840 ();
 sg13g2_fill_2 FILLER_0_149_867 ();
 sg13g2_fill_1 FILLER_0_149_869 ();
 sg13g2_fill_8 FILLER_0_149_896 ();
 sg13g2_fill_8 FILLER_0_149_904 ();
 sg13g2_fill_4 FILLER_0_149_912 ();
 sg13g2_fill_2 FILLER_0_149_916 ();
 sg13g2_fill_8 FILLER_0_149_923 ();
 sg13g2_fill_8 FILLER_0_149_931 ();
 sg13g2_fill_8 FILLER_0_149_939 ();
 sg13g2_fill_8 FILLER_0_149_947 ();
 sg13g2_fill_8 FILLER_0_149_955 ();
 sg13g2_fill_8 FILLER_0_149_963 ();
 sg13g2_fill_8 FILLER_0_149_971 ();
 sg13g2_fill_8 FILLER_0_149_979 ();
 sg13g2_fill_8 FILLER_0_149_987 ();
 sg13g2_fill_1 FILLER_0_149_995 ();
 sg13g2_fill_8 FILLER_0_149_1001 ();
 sg13g2_fill_1 FILLER_0_149_1009 ();
 sg13g2_fill_8 FILLER_0_149_1015 ();
 sg13g2_fill_8 FILLER_0_149_1023 ();
 sg13g2_fill_8 FILLER_0_149_1031 ();
 sg13g2_fill_8 FILLER_0_149_1039 ();
 sg13g2_fill_2 FILLER_0_149_1047 ();
 sg13g2_fill_2 FILLER_0_149_1054 ();
 sg13g2_fill_2 FILLER_0_149_1062 ();
 sg13g2_fill_2 FILLER_0_149_1070 ();
 sg13g2_fill_4 FILLER_0_149_1076 ();
 sg13g2_fill_2 FILLER_0_149_1080 ();
 sg13g2_fill_8 FILLER_0_149_1092 ();
 sg13g2_fill_4 FILLER_0_149_1100 ();
 sg13g2_fill_1 FILLER_0_149_1104 ();
 sg13g2_fill_2 FILLER_0_149_1110 ();
 sg13g2_fill_4 FILLER_0_149_1138 ();
 sg13g2_fill_1 FILLER_0_149_1142 ();
 sg13g2_fill_2 FILLER_0_149_1148 ();
 sg13g2_fill_8 FILLER_0_149_1154 ();
 sg13g2_fill_8 FILLER_0_149_1162 ();
 sg13g2_fill_8 FILLER_0_149_1170 ();
 sg13g2_fill_1 FILLER_0_149_1178 ();
 sg13g2_fill_2 FILLER_0_149_1184 ();
 sg13g2_fill_4 FILLER_0_149_1212 ();
 sg13g2_fill_4 FILLER_0_149_1221 ();
 sg13g2_fill_1 FILLER_0_149_1225 ();
 sg13g2_fill_2 FILLER_0_149_1230 ();
 sg13g2_fill_1 FILLER_0_149_1232 ();
 sg13g2_fill_8 FILLER_0_149_1259 ();
 sg13g2_fill_8 FILLER_0_149_1267 ();
 sg13g2_fill_8 FILLER_0_149_1275 ();
 sg13g2_fill_8 FILLER_0_149_1283 ();
 sg13g2_fill_4 FILLER_0_149_1291 ();
 sg13g2_fill_2 FILLER_0_149_1295 ();
 sg13g2_fill_8 FILLER_0_150_0 ();
 sg13g2_fill_8 FILLER_0_150_8 ();
 sg13g2_fill_8 FILLER_0_150_16 ();
 sg13g2_fill_8 FILLER_0_150_24 ();
 sg13g2_fill_8 FILLER_0_150_32 ();
 sg13g2_fill_8 FILLER_0_150_40 ();
 sg13g2_fill_8 FILLER_0_150_48 ();
 sg13g2_fill_8 FILLER_0_150_56 ();
 sg13g2_fill_8 FILLER_0_150_64 ();
 sg13g2_fill_8 FILLER_0_150_72 ();
 sg13g2_fill_8 FILLER_0_150_80 ();
 sg13g2_fill_8 FILLER_0_150_88 ();
 sg13g2_fill_8 FILLER_0_150_96 ();
 sg13g2_fill_8 FILLER_0_150_104 ();
 sg13g2_fill_8 FILLER_0_150_112 ();
 sg13g2_fill_8 FILLER_0_150_120 ();
 sg13g2_fill_8 FILLER_0_150_128 ();
 sg13g2_fill_8 FILLER_0_150_136 ();
 sg13g2_fill_8 FILLER_0_150_144 ();
 sg13g2_fill_8 FILLER_0_150_152 ();
 sg13g2_fill_8 FILLER_0_150_160 ();
 sg13g2_fill_8 FILLER_0_150_168 ();
 sg13g2_fill_8 FILLER_0_150_176 ();
 sg13g2_fill_8 FILLER_0_150_184 ();
 sg13g2_fill_8 FILLER_0_150_192 ();
 sg13g2_fill_8 FILLER_0_150_200 ();
 sg13g2_fill_8 FILLER_0_150_208 ();
 sg13g2_fill_8 FILLER_0_150_216 ();
 sg13g2_fill_8 FILLER_0_150_224 ();
 sg13g2_fill_8 FILLER_0_150_232 ();
 sg13g2_fill_8 FILLER_0_150_240 ();
 sg13g2_fill_8 FILLER_0_150_248 ();
 sg13g2_fill_8 FILLER_0_150_256 ();
 sg13g2_fill_8 FILLER_0_150_264 ();
 sg13g2_fill_8 FILLER_0_150_272 ();
 sg13g2_fill_8 FILLER_0_150_280 ();
 sg13g2_fill_8 FILLER_0_150_288 ();
 sg13g2_fill_1 FILLER_0_150_296 ();
 sg13g2_fill_8 FILLER_0_150_302 ();
 sg13g2_fill_1 FILLER_0_150_310 ();
 sg13g2_fill_8 FILLER_0_150_315 ();
 sg13g2_fill_4 FILLER_0_150_323 ();
 sg13g2_fill_8 FILLER_0_150_353 ();
 sg13g2_fill_4 FILLER_0_150_361 ();
 sg13g2_fill_1 FILLER_0_150_365 ();
 sg13g2_fill_8 FILLER_0_150_370 ();
 sg13g2_fill_8 FILLER_0_150_378 ();
 sg13g2_fill_4 FILLER_0_150_386 ();
 sg13g2_fill_2 FILLER_0_150_390 ();
 sg13g2_fill_4 FILLER_0_150_396 ();
 sg13g2_fill_1 FILLER_0_150_400 ();
 sg13g2_fill_2 FILLER_0_150_406 ();
 sg13g2_fill_4 FILLER_0_150_412 ();
 sg13g2_fill_2 FILLER_0_150_416 ();
 sg13g2_fill_4 FILLER_0_150_444 ();
 sg13g2_fill_2 FILLER_0_150_448 ();
 sg13g2_fill_8 FILLER_0_150_455 ();
 sg13g2_fill_8 FILLER_0_150_468 ();
 sg13g2_fill_4 FILLER_0_150_476 ();
 sg13g2_fill_8 FILLER_0_150_501 ();
 sg13g2_fill_4 FILLER_0_150_509 ();
 sg13g2_fill_1 FILLER_0_150_513 ();
 sg13g2_fill_2 FILLER_0_150_518 ();
 sg13g2_fill_4 FILLER_0_150_546 ();
 sg13g2_fill_2 FILLER_0_150_550 ();
 sg13g2_fill_1 FILLER_0_150_552 ();
 sg13g2_fill_8 FILLER_0_150_579 ();
 sg13g2_fill_2 FILLER_0_150_587 ();
 sg13g2_fill_1 FILLER_0_150_589 ();
 sg13g2_fill_4 FILLER_0_150_595 ();
 sg13g2_fill_4 FILLER_0_150_604 ();
 sg13g2_fill_4 FILLER_0_150_613 ();
 sg13g2_fill_2 FILLER_0_150_622 ();
 sg13g2_fill_8 FILLER_0_150_628 ();
 sg13g2_fill_8 FILLER_0_150_636 ();
 sg13g2_fill_8 FILLER_0_150_649 ();
 sg13g2_fill_8 FILLER_0_150_657 ();
 sg13g2_fill_2 FILLER_0_150_665 ();
 sg13g2_fill_8 FILLER_0_150_679 ();
 sg13g2_fill_8 FILLER_0_150_687 ();
 sg13g2_fill_2 FILLER_0_150_695 ();
 sg13g2_fill_8 FILLER_0_150_702 ();
 sg13g2_fill_8 FILLER_0_150_710 ();
 sg13g2_fill_8 FILLER_0_150_718 ();
 sg13g2_fill_4 FILLER_0_150_731 ();
 sg13g2_fill_2 FILLER_0_150_739 ();
 sg13g2_fill_2 FILLER_0_150_767 ();
 sg13g2_fill_8 FILLER_0_150_773 ();
 sg13g2_fill_8 FILLER_0_150_781 ();
 sg13g2_fill_4 FILLER_0_150_789 ();
 sg13g2_fill_2 FILLER_0_150_798 ();
 sg13g2_fill_8 FILLER_0_150_804 ();
 sg13g2_fill_2 FILLER_0_150_817 ();
 sg13g2_fill_4 FILLER_0_150_824 ();
 sg13g2_fill_1 FILLER_0_150_828 ();
 sg13g2_fill_2 FILLER_0_150_834 ();
 sg13g2_fill_4 FILLER_0_150_862 ();
 sg13g2_fill_8 FILLER_0_150_887 ();
 sg13g2_fill_8 FILLER_0_150_895 ();
 sg13g2_fill_4 FILLER_0_150_903 ();
 sg13g2_fill_1 FILLER_0_150_907 ();
 sg13g2_fill_2 FILLER_0_150_913 ();
 sg13g2_fill_8 FILLER_0_150_920 ();
 sg13g2_fill_8 FILLER_0_150_928 ();
 sg13g2_fill_4 FILLER_0_150_936 ();
 sg13g2_fill_2 FILLER_0_150_944 ();
 sg13g2_fill_8 FILLER_0_150_972 ();
 sg13g2_fill_2 FILLER_0_150_980 ();
 sg13g2_fill_1 FILLER_0_150_982 ();
 sg13g2_fill_2 FILLER_0_150_988 ();
 sg13g2_fill_1 FILLER_0_150_990 ();
 sg13g2_fill_2 FILLER_0_150_996 ();
 sg13g2_fill_1 FILLER_0_150_998 ();
 sg13g2_fill_2 FILLER_0_150_1005 ();
 sg13g2_fill_8 FILLER_0_150_1011 ();
 sg13g2_fill_4 FILLER_0_150_1019 ();
 sg13g2_fill_1 FILLER_0_150_1023 ();
 sg13g2_fill_8 FILLER_0_150_1029 ();
 sg13g2_fill_8 FILLER_0_150_1037 ();
 sg13g2_fill_8 FILLER_0_150_1045 ();
 sg13g2_fill_4 FILLER_0_150_1053 ();
 sg13g2_fill_2 FILLER_0_150_1062 ();
 sg13g2_fill_2 FILLER_0_150_1090 ();
 sg13g2_fill_4 FILLER_0_150_1097 ();
 sg13g2_fill_2 FILLER_0_150_1106 ();
 sg13g2_fill_2 FILLER_0_150_1112 ();
 sg13g2_fill_2 FILLER_0_150_1140 ();
 sg13g2_fill_8 FILLER_0_150_1168 ();
 sg13g2_fill_4 FILLER_0_150_1176 ();
 sg13g2_fill_1 FILLER_0_150_1180 ();
 sg13g2_fill_8 FILLER_0_150_1186 ();
 sg13g2_fill_8 FILLER_0_150_1194 ();
 sg13g2_fill_8 FILLER_0_150_1202 ();
 sg13g2_fill_2 FILLER_0_150_1210 ();
 sg13g2_fill_8 FILLER_0_150_1217 ();
 sg13g2_fill_4 FILLER_0_150_1225 ();
 sg13g2_fill_2 FILLER_0_150_1229 ();
 sg13g2_fill_2 FILLER_0_150_1236 ();
 sg13g2_fill_8 FILLER_0_150_1242 ();
 sg13g2_fill_8 FILLER_0_150_1250 ();
 sg13g2_fill_8 FILLER_0_150_1258 ();
 sg13g2_fill_8 FILLER_0_150_1266 ();
 sg13g2_fill_8 FILLER_0_150_1274 ();
 sg13g2_fill_8 FILLER_0_150_1282 ();
 sg13g2_fill_4 FILLER_0_150_1290 ();
 sg13g2_fill_2 FILLER_0_150_1294 ();
 sg13g2_fill_1 FILLER_0_150_1296 ();
 sg13g2_fill_8 FILLER_0_151_0 ();
 sg13g2_fill_8 FILLER_0_151_8 ();
 sg13g2_fill_8 FILLER_0_151_16 ();
 sg13g2_fill_8 FILLER_0_151_24 ();
 sg13g2_fill_8 FILLER_0_151_32 ();
 sg13g2_fill_8 FILLER_0_151_40 ();
 sg13g2_fill_8 FILLER_0_151_48 ();
 sg13g2_fill_8 FILLER_0_151_56 ();
 sg13g2_fill_8 FILLER_0_151_64 ();
 sg13g2_fill_8 FILLER_0_151_72 ();
 sg13g2_fill_8 FILLER_0_151_80 ();
 sg13g2_fill_8 FILLER_0_151_88 ();
 sg13g2_fill_8 FILLER_0_151_96 ();
 sg13g2_fill_8 FILLER_0_151_104 ();
 sg13g2_fill_8 FILLER_0_151_112 ();
 sg13g2_fill_8 FILLER_0_151_120 ();
 sg13g2_fill_8 FILLER_0_151_128 ();
 sg13g2_fill_8 FILLER_0_151_136 ();
 sg13g2_fill_8 FILLER_0_151_144 ();
 sg13g2_fill_8 FILLER_0_151_152 ();
 sg13g2_fill_8 FILLER_0_151_160 ();
 sg13g2_fill_8 FILLER_0_151_168 ();
 sg13g2_fill_8 FILLER_0_151_176 ();
 sg13g2_fill_8 FILLER_0_151_184 ();
 sg13g2_fill_8 FILLER_0_151_192 ();
 sg13g2_fill_8 FILLER_0_151_200 ();
 sg13g2_fill_8 FILLER_0_151_208 ();
 sg13g2_fill_8 FILLER_0_151_216 ();
 sg13g2_fill_8 FILLER_0_151_224 ();
 sg13g2_fill_8 FILLER_0_151_232 ();
 sg13g2_fill_8 FILLER_0_151_240 ();
 sg13g2_fill_8 FILLER_0_151_248 ();
 sg13g2_fill_8 FILLER_0_151_256 ();
 sg13g2_fill_8 FILLER_0_151_264 ();
 sg13g2_fill_8 FILLER_0_151_272 ();
 sg13g2_fill_4 FILLER_0_151_280 ();
 sg13g2_fill_2 FILLER_0_151_284 ();
 sg13g2_fill_2 FILLER_0_151_291 ();
 sg13g2_fill_2 FILLER_0_151_319 ();
 sg13g2_fill_1 FILLER_0_151_321 ();
 sg13g2_fill_8 FILLER_0_151_327 ();
 sg13g2_fill_4 FILLER_0_151_335 ();
 sg13g2_fill_2 FILLER_0_151_344 ();
 sg13g2_fill_8 FILLER_0_151_350 ();
 sg13g2_fill_4 FILLER_0_151_358 ();
 sg13g2_fill_2 FILLER_0_151_362 ();
 sg13g2_fill_8 FILLER_0_151_369 ();
 sg13g2_fill_4 FILLER_0_151_377 ();
 sg13g2_fill_2 FILLER_0_151_381 ();
 sg13g2_fill_8 FILLER_0_151_388 ();
 sg13g2_fill_4 FILLER_0_151_396 ();
 sg13g2_fill_2 FILLER_0_151_426 ();
 sg13g2_fill_2 FILLER_0_151_449 ();
 sg13g2_fill_8 FILLER_0_151_456 ();
 sg13g2_fill_2 FILLER_0_151_464 ();
 sg13g2_fill_1 FILLER_0_151_466 ();
 sg13g2_fill_8 FILLER_0_151_493 ();
 sg13g2_fill_4 FILLER_0_151_501 ();
 sg13g2_fill_1 FILLER_0_151_505 ();
 sg13g2_fill_2 FILLER_0_151_511 ();
 sg13g2_fill_2 FILLER_0_151_539 ();
 sg13g2_fill_1 FILLER_0_151_541 ();
 sg13g2_fill_4 FILLER_0_151_547 ();
 sg13g2_fill_8 FILLER_0_151_555 ();
 sg13g2_fill_8 FILLER_0_151_563 ();
 sg13g2_fill_8 FILLER_0_151_571 ();
 sg13g2_fill_8 FILLER_0_151_579 ();
 sg13g2_fill_8 FILLER_0_151_587 ();
 sg13g2_fill_8 FILLER_0_151_595 ();
 sg13g2_fill_8 FILLER_0_151_603 ();
 sg13g2_fill_8 FILLER_0_151_611 ();
 sg13g2_fill_8 FILLER_0_151_619 ();
 sg13g2_fill_8 FILLER_0_151_627 ();
 sg13g2_fill_1 FILLER_0_151_635 ();
 sg13g2_fill_2 FILLER_0_151_641 ();
 sg13g2_fill_8 FILLER_0_151_648 ();
 sg13g2_fill_8 FILLER_0_151_656 ();
 sg13g2_fill_8 FILLER_0_151_664 ();
 sg13g2_fill_4 FILLER_0_151_672 ();
 sg13g2_fill_2 FILLER_0_151_676 ();
 sg13g2_fill_2 FILLER_0_151_683 ();
 sg13g2_fill_8 FILLER_0_151_689 ();
 sg13g2_fill_8 FILLER_0_151_697 ();
 sg13g2_fill_8 FILLER_0_151_705 ();
 sg13g2_fill_4 FILLER_0_151_713 ();
 sg13g2_fill_1 FILLER_0_151_717 ();
 sg13g2_fill_8 FILLER_0_151_744 ();
 sg13g2_fill_8 FILLER_0_151_773 ();
 sg13g2_fill_8 FILLER_0_151_781 ();
 sg13g2_fill_8 FILLER_0_151_789 ();
 sg13g2_fill_8 FILLER_0_151_797 ();
 sg13g2_fill_4 FILLER_0_151_805 ();
 sg13g2_fill_2 FILLER_0_151_809 ();
 sg13g2_fill_8 FILLER_0_151_816 ();
 sg13g2_fill_8 FILLER_0_151_824 ();
 sg13g2_fill_1 FILLER_0_151_832 ();
 sg13g2_fill_2 FILLER_0_151_837 ();
 sg13g2_fill_2 FILLER_0_151_844 ();
 sg13g2_fill_2 FILLER_0_151_850 ();
 sg13g2_fill_2 FILLER_0_151_878 ();
 sg13g2_fill_8 FILLER_0_151_887 ();
 sg13g2_fill_2 FILLER_0_151_900 ();
 sg13g2_fill_2 FILLER_0_151_928 ();
 sg13g2_fill_4 FILLER_0_151_935 ();
 sg13g2_fill_2 FILLER_0_151_939 ();
 sg13g2_fill_1 FILLER_0_151_941 ();
 sg13g2_fill_2 FILLER_0_151_947 ();
 sg13g2_fill_2 FILLER_0_151_975 ();
 sg13g2_fill_4 FILLER_0_151_982 ();
 sg13g2_fill_4 FILLER_0_151_1012 ();
 sg13g2_fill_2 FILLER_0_151_1021 ();
 sg13g2_fill_1 FILLER_0_151_1023 ();
 sg13g2_fill_2 FILLER_0_151_1029 ();
 sg13g2_fill_8 FILLER_0_151_1039 ();
 sg13g2_fill_8 FILLER_0_151_1047 ();
 sg13g2_fill_2 FILLER_0_151_1055 ();
 sg13g2_fill_2 FILLER_0_151_1062 ();
 sg13g2_fill_8 FILLER_0_151_1069 ();
 sg13g2_fill_8 FILLER_0_151_1077 ();
 sg13g2_fill_8 FILLER_0_151_1085 ();
 sg13g2_fill_4 FILLER_0_151_1093 ();
 sg13g2_fill_2 FILLER_0_151_1097 ();
 sg13g2_fill_1 FILLER_0_151_1099 ();
 sg13g2_fill_2 FILLER_0_151_1106 ();
 sg13g2_fill_4 FILLER_0_151_1113 ();
 sg13g2_fill_1 FILLER_0_151_1117 ();
 sg13g2_fill_4 FILLER_0_151_1123 ();
 sg13g2_fill_8 FILLER_0_151_1131 ();
 sg13g2_fill_2 FILLER_0_151_1160 ();
 sg13g2_fill_8 FILLER_0_151_1168 ();
 sg13g2_fill_8 FILLER_0_151_1176 ();
 sg13g2_fill_8 FILLER_0_151_1184 ();
 sg13g2_fill_8 FILLER_0_151_1192 ();
 sg13g2_fill_8 FILLER_0_151_1200 ();
 sg13g2_fill_8 FILLER_0_151_1208 ();
 sg13g2_fill_8 FILLER_0_151_1216 ();
 sg13g2_fill_8 FILLER_0_151_1224 ();
 sg13g2_fill_8 FILLER_0_151_1232 ();
 sg13g2_fill_8 FILLER_0_151_1240 ();
 sg13g2_fill_8 FILLER_0_151_1248 ();
 sg13g2_fill_8 FILLER_0_151_1256 ();
 sg13g2_fill_8 FILLER_0_151_1264 ();
 sg13g2_fill_8 FILLER_0_151_1272 ();
 sg13g2_fill_8 FILLER_0_151_1280 ();
 sg13g2_fill_8 FILLER_0_151_1288 ();
 sg13g2_fill_1 FILLER_0_151_1296 ();
 sg13g2_fill_8 FILLER_0_152_0 ();
 sg13g2_fill_8 FILLER_0_152_8 ();
 sg13g2_fill_8 FILLER_0_152_16 ();
 sg13g2_fill_8 FILLER_0_152_24 ();
 sg13g2_fill_8 FILLER_0_152_32 ();
 sg13g2_fill_8 FILLER_0_152_40 ();
 sg13g2_fill_8 FILLER_0_152_48 ();
 sg13g2_fill_8 FILLER_0_152_56 ();
 sg13g2_fill_8 FILLER_0_152_64 ();
 sg13g2_fill_8 FILLER_0_152_72 ();
 sg13g2_fill_8 FILLER_0_152_80 ();
 sg13g2_fill_8 FILLER_0_152_88 ();
 sg13g2_fill_8 FILLER_0_152_96 ();
 sg13g2_fill_8 FILLER_0_152_104 ();
 sg13g2_fill_8 FILLER_0_152_112 ();
 sg13g2_fill_8 FILLER_0_152_120 ();
 sg13g2_fill_8 FILLER_0_152_128 ();
 sg13g2_fill_8 FILLER_0_152_136 ();
 sg13g2_fill_8 FILLER_0_152_144 ();
 sg13g2_fill_8 FILLER_0_152_152 ();
 sg13g2_fill_8 FILLER_0_152_160 ();
 sg13g2_fill_8 FILLER_0_152_168 ();
 sg13g2_fill_8 FILLER_0_152_176 ();
 sg13g2_fill_8 FILLER_0_152_184 ();
 sg13g2_fill_8 FILLER_0_152_192 ();
 sg13g2_fill_8 FILLER_0_152_200 ();
 sg13g2_fill_8 FILLER_0_152_208 ();
 sg13g2_fill_8 FILLER_0_152_216 ();
 sg13g2_fill_8 FILLER_0_152_224 ();
 sg13g2_fill_8 FILLER_0_152_232 ();
 sg13g2_fill_8 FILLER_0_152_240 ();
 sg13g2_fill_8 FILLER_0_152_248 ();
 sg13g2_fill_8 FILLER_0_152_256 ();
 sg13g2_fill_8 FILLER_0_152_264 ();
 sg13g2_fill_8 FILLER_0_152_272 ();
 sg13g2_fill_8 FILLER_0_152_280 ();
 sg13g2_fill_8 FILLER_0_152_288 ();
 sg13g2_fill_8 FILLER_0_152_296 ();
 sg13g2_fill_8 FILLER_0_152_304 ();
 sg13g2_fill_4 FILLER_0_152_312 ();
 sg13g2_fill_1 FILLER_0_152_316 ();
 sg13g2_fill_8 FILLER_0_152_320 ();
 sg13g2_fill_8 FILLER_0_152_328 ();
 sg13g2_fill_8 FILLER_0_152_362 ();
 sg13g2_fill_4 FILLER_0_152_370 ();
 sg13g2_fill_1 FILLER_0_152_374 ();
 sg13g2_fill_2 FILLER_0_152_401 ();
 sg13g2_fill_4 FILLER_0_152_408 ();
 sg13g2_fill_2 FILLER_0_152_412 ();
 sg13g2_fill_1 FILLER_0_152_414 ();
 sg13g2_fill_4 FILLER_0_152_421 ();
 sg13g2_fill_1 FILLER_0_152_425 ();
 sg13g2_fill_4 FILLER_0_152_431 ();
 sg13g2_fill_2 FILLER_0_152_440 ();
 sg13g2_fill_8 FILLER_0_152_447 ();
 sg13g2_fill_8 FILLER_0_152_455 ();
 sg13g2_fill_2 FILLER_0_152_463 ();
 sg13g2_fill_8 FILLER_0_152_491 ();
 sg13g2_fill_8 FILLER_0_152_499 ();
 sg13g2_fill_8 FILLER_0_152_507 ();
 sg13g2_fill_8 FILLER_0_152_515 ();
 sg13g2_fill_8 FILLER_0_152_523 ();
 sg13g2_fill_1 FILLER_0_152_531 ();
 sg13g2_fill_2 FILLER_0_152_558 ();
 sg13g2_fill_4 FILLER_0_152_565 ();
 sg13g2_fill_2 FILLER_0_152_569 ();
 sg13g2_fill_8 FILLER_0_152_581 ();
 sg13g2_fill_8 FILLER_0_152_589 ();
 sg13g2_fill_8 FILLER_0_152_597 ();
 sg13g2_fill_8 FILLER_0_152_605 ();
 sg13g2_fill_8 FILLER_0_152_613 ();
 sg13g2_fill_4 FILLER_0_152_621 ();
 sg13g2_fill_2 FILLER_0_152_625 ();
 sg13g2_fill_1 FILLER_0_152_627 ();
 sg13g2_fill_4 FILLER_0_152_638 ();
 sg13g2_fill_2 FILLER_0_152_642 ();
 sg13g2_fill_8 FILLER_0_152_650 ();
 sg13g2_fill_4 FILLER_0_152_658 ();
 sg13g2_fill_1 FILLER_0_152_662 ();
 sg13g2_fill_4 FILLER_0_152_668 ();
 sg13g2_fill_1 FILLER_0_152_672 ();
 sg13g2_fill_2 FILLER_0_152_679 ();
 sg13g2_fill_8 FILLER_0_152_707 ();
 sg13g2_fill_2 FILLER_0_152_715 ();
 sg13g2_fill_4 FILLER_0_152_743 ();
 sg13g2_fill_4 FILLER_0_152_768 ();
 sg13g2_fill_1 FILLER_0_152_772 ();
 sg13g2_fill_4 FILLER_0_152_779 ();
 sg13g2_fill_1 FILLER_0_152_783 ();
 sg13g2_fill_4 FILLER_0_152_788 ();
 sg13g2_fill_8 FILLER_0_152_796 ();
 sg13g2_fill_8 FILLER_0_152_804 ();
 sg13g2_fill_8 FILLER_0_152_812 ();
 sg13g2_fill_8 FILLER_0_152_820 ();
 sg13g2_fill_8 FILLER_0_152_828 ();
 sg13g2_fill_8 FILLER_0_152_841 ();
 sg13g2_fill_8 FILLER_0_152_849 ();
 sg13g2_fill_8 FILLER_0_152_857 ();
 sg13g2_fill_8 FILLER_0_152_865 ();
 sg13g2_fill_4 FILLER_0_152_878 ();
 sg13g2_fill_8 FILLER_0_152_886 ();
 sg13g2_fill_8 FILLER_0_152_894 ();
 sg13g2_fill_8 FILLER_0_152_902 ();
 sg13g2_fill_1 FILLER_0_152_910 ();
 sg13g2_fill_8 FILLER_0_152_916 ();
 sg13g2_fill_1 FILLER_0_152_924 ();
 sg13g2_fill_8 FILLER_0_152_929 ();
 sg13g2_fill_4 FILLER_0_152_937 ();
 sg13g2_fill_1 FILLER_0_152_941 ();
 sg13g2_fill_2 FILLER_0_152_949 ();
 sg13g2_fill_2 FILLER_0_152_956 ();
 sg13g2_fill_2 FILLER_0_152_962 ();
 sg13g2_fill_1 FILLER_0_152_964 ();
 sg13g2_fill_4 FILLER_0_152_975 ();
 sg13g2_fill_8 FILLER_0_152_984 ();
 sg13g2_fill_4 FILLER_0_152_992 ();
 sg13g2_fill_2 FILLER_0_152_996 ();
 sg13g2_fill_2 FILLER_0_152_1004 ();
 sg13g2_fill_8 FILLER_0_152_1011 ();
 sg13g2_fill_8 FILLER_0_152_1019 ();
 sg13g2_fill_8 FILLER_0_152_1033 ();
 sg13g2_fill_8 FILLER_0_152_1041 ();
 sg13g2_fill_8 FILLER_0_152_1049 ();
 sg13g2_fill_2 FILLER_0_152_1057 ();
 sg13g2_fill_1 FILLER_0_152_1059 ();
 sg13g2_fill_8 FILLER_0_152_1086 ();
 sg13g2_fill_8 FILLER_0_152_1094 ();
 sg13g2_fill_8 FILLER_0_152_1102 ();
 sg13g2_fill_2 FILLER_0_152_1110 ();
 sg13g2_fill_2 FILLER_0_152_1120 ();
 sg13g2_fill_2 FILLER_0_152_1127 ();
 sg13g2_fill_2 FILLER_0_152_1155 ();
 sg13g2_fill_1 FILLER_0_152_1157 ();
 sg13g2_fill_2 FILLER_0_152_1162 ();
 sg13g2_fill_2 FILLER_0_152_1169 ();
 sg13g2_fill_1 FILLER_0_152_1171 ();
 sg13g2_fill_2 FILLER_0_152_1176 ();
 sg13g2_fill_2 FILLER_0_152_1183 ();
 sg13g2_fill_8 FILLER_0_152_1211 ();
 sg13g2_fill_8 FILLER_0_152_1219 ();
 sg13g2_fill_8 FILLER_0_152_1227 ();
 sg13g2_fill_8 FILLER_0_152_1235 ();
 sg13g2_fill_8 FILLER_0_152_1243 ();
 sg13g2_fill_8 FILLER_0_152_1251 ();
 sg13g2_fill_8 FILLER_0_152_1259 ();
 sg13g2_fill_8 FILLER_0_152_1267 ();
 sg13g2_fill_8 FILLER_0_152_1275 ();
 sg13g2_fill_8 FILLER_0_152_1283 ();
 sg13g2_fill_4 FILLER_0_152_1291 ();
 sg13g2_fill_2 FILLER_0_152_1295 ();
 sg13g2_fill_8 FILLER_0_153_0 ();
 sg13g2_fill_8 FILLER_0_153_8 ();
 sg13g2_fill_8 FILLER_0_153_16 ();
 sg13g2_fill_8 FILLER_0_153_24 ();
 sg13g2_fill_8 FILLER_0_153_32 ();
 sg13g2_fill_8 FILLER_0_153_40 ();
 sg13g2_fill_8 FILLER_0_153_48 ();
 sg13g2_fill_8 FILLER_0_153_56 ();
 sg13g2_fill_8 FILLER_0_153_64 ();
 sg13g2_fill_8 FILLER_0_153_72 ();
 sg13g2_fill_8 FILLER_0_153_80 ();
 sg13g2_fill_8 FILLER_0_153_88 ();
 sg13g2_fill_8 FILLER_0_153_96 ();
 sg13g2_fill_8 FILLER_0_153_104 ();
 sg13g2_fill_8 FILLER_0_153_112 ();
 sg13g2_fill_8 FILLER_0_153_120 ();
 sg13g2_fill_8 FILLER_0_153_128 ();
 sg13g2_fill_8 FILLER_0_153_136 ();
 sg13g2_fill_8 FILLER_0_153_144 ();
 sg13g2_fill_8 FILLER_0_153_152 ();
 sg13g2_fill_8 FILLER_0_153_160 ();
 sg13g2_fill_8 FILLER_0_153_168 ();
 sg13g2_fill_8 FILLER_0_153_176 ();
 sg13g2_fill_8 FILLER_0_153_184 ();
 sg13g2_fill_8 FILLER_0_153_192 ();
 sg13g2_fill_8 FILLER_0_153_200 ();
 sg13g2_fill_8 FILLER_0_153_208 ();
 sg13g2_fill_8 FILLER_0_153_216 ();
 sg13g2_fill_8 FILLER_0_153_224 ();
 sg13g2_fill_8 FILLER_0_153_232 ();
 sg13g2_fill_8 FILLER_0_153_240 ();
 sg13g2_fill_8 FILLER_0_153_248 ();
 sg13g2_fill_8 FILLER_0_153_256 ();
 sg13g2_fill_8 FILLER_0_153_264 ();
 sg13g2_fill_8 FILLER_0_153_272 ();
 sg13g2_fill_8 FILLER_0_153_280 ();
 sg13g2_fill_8 FILLER_0_153_288 ();
 sg13g2_fill_8 FILLER_0_153_296 ();
 sg13g2_fill_8 FILLER_0_153_304 ();
 sg13g2_fill_8 FILLER_0_153_312 ();
 sg13g2_fill_8 FILLER_0_153_320 ();
 sg13g2_fill_8 FILLER_0_153_328 ();
 sg13g2_fill_8 FILLER_0_153_336 ();
 sg13g2_fill_8 FILLER_0_153_344 ();
 sg13g2_fill_2 FILLER_0_153_373 ();
 sg13g2_fill_2 FILLER_0_153_385 ();
 sg13g2_fill_4 FILLER_0_153_391 ();
 sg13g2_fill_1 FILLER_0_153_395 ();
 sg13g2_fill_2 FILLER_0_153_401 ();
 sg13g2_fill_8 FILLER_0_153_409 ();
 sg13g2_fill_8 FILLER_0_153_417 ();
 sg13g2_fill_8 FILLER_0_153_425 ();
 sg13g2_fill_8 FILLER_0_153_433 ();
 sg13g2_fill_8 FILLER_0_153_441 ();
 sg13g2_fill_8 FILLER_0_153_449 ();
 sg13g2_fill_2 FILLER_0_153_457 ();
 sg13g2_fill_1 FILLER_0_153_459 ();
 sg13g2_fill_2 FILLER_0_153_465 ();
 sg13g2_fill_4 FILLER_0_153_472 ();
 sg13g2_fill_2 FILLER_0_153_480 ();
 sg13g2_fill_1 FILLER_0_153_482 ();
 sg13g2_fill_8 FILLER_0_153_487 ();
 sg13g2_fill_4 FILLER_0_153_495 ();
 sg13g2_fill_1 FILLER_0_153_499 ();
 sg13g2_fill_8 FILLER_0_153_505 ();
 sg13g2_fill_1 FILLER_0_153_513 ();
 sg13g2_fill_8 FILLER_0_153_518 ();
 sg13g2_fill_2 FILLER_0_153_526 ();
 sg13g2_fill_4 FILLER_0_153_549 ();
 sg13g2_fill_2 FILLER_0_153_553 ();
 sg13g2_fill_1 FILLER_0_153_555 ();
 sg13g2_fill_2 FILLER_0_153_577 ();
 sg13g2_fill_8 FILLER_0_153_583 ();
 sg13g2_fill_8 FILLER_0_153_591 ();
 sg13g2_fill_4 FILLER_0_153_599 ();
 sg13g2_fill_2 FILLER_0_153_603 ();
 sg13g2_fill_2 FILLER_0_153_610 ();
 sg13g2_fill_1 FILLER_0_153_612 ();
 sg13g2_fill_2 FILLER_0_153_639 ();
 sg13g2_fill_2 FILLER_0_153_647 ();
 sg13g2_fill_2 FILLER_0_153_655 ();
 sg13g2_fill_4 FILLER_0_153_661 ();
 sg13g2_fill_1 FILLER_0_153_665 ();
 sg13g2_fill_2 FILLER_0_153_692 ();
 sg13g2_fill_8 FILLER_0_153_698 ();
 sg13g2_fill_8 FILLER_0_153_706 ();
 sg13g2_fill_8 FILLER_0_153_714 ();
 sg13g2_fill_4 FILLER_0_153_722 ();
 sg13g2_fill_2 FILLER_0_153_731 ();
 sg13g2_fill_1 FILLER_0_153_733 ();
 sg13g2_fill_8 FILLER_0_153_738 ();
 sg13g2_fill_8 FILLER_0_153_746 ();
 sg13g2_fill_8 FILLER_0_153_754 ();
 sg13g2_fill_8 FILLER_0_153_762 ();
 sg13g2_fill_8 FILLER_0_153_770 ();
 sg13g2_fill_8 FILLER_0_153_783 ();
 sg13g2_fill_1 FILLER_0_153_791 ();
 sg13g2_fill_2 FILLER_0_153_797 ();
 sg13g2_fill_2 FILLER_0_153_805 ();
 sg13g2_fill_2 FILLER_0_153_814 ();
 sg13g2_fill_8 FILLER_0_153_821 ();
 sg13g2_fill_8 FILLER_0_153_829 ();
 sg13g2_fill_8 FILLER_0_153_837 ();
 sg13g2_fill_8 FILLER_0_153_845 ();
 sg13g2_fill_8 FILLER_0_153_853 ();
 sg13g2_fill_8 FILLER_0_153_861 ();
 sg13g2_fill_8 FILLER_0_153_869 ();
 sg13g2_fill_2 FILLER_0_153_877 ();
 sg13g2_fill_4 FILLER_0_153_884 ();
 sg13g2_fill_2 FILLER_0_153_896 ();
 sg13g2_fill_2 FILLER_0_153_903 ();
 sg13g2_fill_1 FILLER_0_153_905 ();
 sg13g2_fill_8 FILLER_0_153_912 ();
 sg13g2_fill_8 FILLER_0_153_920 ();
 sg13g2_fill_8 FILLER_0_153_928 ();
 sg13g2_fill_8 FILLER_0_153_936 ();
 sg13g2_fill_8 FILLER_0_153_944 ();
 sg13g2_fill_8 FILLER_0_153_952 ();
 sg13g2_fill_8 FILLER_0_153_960 ();
 sg13g2_fill_8 FILLER_0_153_968 ();
 sg13g2_fill_4 FILLER_0_153_976 ();
 sg13g2_fill_2 FILLER_0_153_980 ();
 sg13g2_fill_8 FILLER_0_153_987 ();
 sg13g2_fill_8 FILLER_0_153_995 ();
 sg13g2_fill_8 FILLER_0_153_1003 ();
 sg13g2_fill_8 FILLER_0_153_1011 ();
 sg13g2_fill_8 FILLER_0_153_1019 ();
 sg13g2_fill_2 FILLER_0_153_1032 ();
 sg13g2_fill_8 FILLER_0_153_1038 ();
 sg13g2_fill_8 FILLER_0_153_1046 ();
 sg13g2_fill_4 FILLER_0_153_1054 ();
 sg13g2_fill_2 FILLER_0_153_1058 ();
 sg13g2_fill_1 FILLER_0_153_1060 ();
 sg13g2_fill_2 FILLER_0_153_1066 ();
 sg13g2_fill_8 FILLER_0_153_1072 ();
 sg13g2_fill_8 FILLER_0_153_1080 ();
 sg13g2_fill_8 FILLER_0_153_1088 ();
 sg13g2_fill_8 FILLER_0_153_1096 ();
 sg13g2_fill_8 FILLER_0_153_1104 ();
 sg13g2_fill_8 FILLER_0_153_1112 ();
 sg13g2_fill_8 FILLER_0_153_1120 ();
 sg13g2_fill_8 FILLER_0_153_1128 ();
 sg13g2_fill_8 FILLER_0_153_1136 ();
 sg13g2_fill_8 FILLER_0_153_1144 ();
 sg13g2_fill_8 FILLER_0_153_1152 ();
 sg13g2_fill_8 FILLER_0_153_1160 ();
 sg13g2_fill_8 FILLER_0_153_1168 ();
 sg13g2_fill_4 FILLER_0_153_1176 ();
 sg13g2_fill_1 FILLER_0_153_1180 ();
 sg13g2_fill_2 FILLER_0_153_1186 ();
 sg13g2_fill_8 FILLER_0_153_1214 ();
 sg13g2_fill_2 FILLER_0_153_1222 ();
 sg13g2_fill_1 FILLER_0_153_1224 ();
 sg13g2_fill_2 FILLER_0_153_1229 ();
 sg13g2_fill_8 FILLER_0_153_1257 ();
 sg13g2_fill_8 FILLER_0_153_1265 ();
 sg13g2_fill_8 FILLER_0_153_1273 ();
 sg13g2_fill_8 FILLER_0_153_1281 ();
 sg13g2_fill_8 FILLER_0_153_1289 ();
 sg13g2_fill_8 FILLER_0_154_0 ();
 sg13g2_fill_8 FILLER_0_154_8 ();
 sg13g2_fill_8 FILLER_0_154_16 ();
 sg13g2_fill_8 FILLER_0_154_24 ();
 sg13g2_fill_8 FILLER_0_154_32 ();
 sg13g2_fill_8 FILLER_0_154_40 ();
 sg13g2_fill_8 FILLER_0_154_48 ();
 sg13g2_fill_8 FILLER_0_154_56 ();
 sg13g2_fill_8 FILLER_0_154_64 ();
 sg13g2_fill_8 FILLER_0_154_72 ();
 sg13g2_fill_8 FILLER_0_154_80 ();
 sg13g2_fill_8 FILLER_0_154_88 ();
 sg13g2_fill_8 FILLER_0_154_96 ();
 sg13g2_fill_8 FILLER_0_154_104 ();
 sg13g2_fill_8 FILLER_0_154_112 ();
 sg13g2_fill_8 FILLER_0_154_120 ();
 sg13g2_fill_8 FILLER_0_154_128 ();
 sg13g2_fill_8 FILLER_0_154_136 ();
 sg13g2_fill_8 FILLER_0_154_144 ();
 sg13g2_fill_8 FILLER_0_154_152 ();
 sg13g2_fill_8 FILLER_0_154_160 ();
 sg13g2_fill_8 FILLER_0_154_168 ();
 sg13g2_fill_8 FILLER_0_154_176 ();
 sg13g2_fill_8 FILLER_0_154_184 ();
 sg13g2_fill_8 FILLER_0_154_192 ();
 sg13g2_fill_8 FILLER_0_154_200 ();
 sg13g2_fill_8 FILLER_0_154_208 ();
 sg13g2_fill_8 FILLER_0_154_216 ();
 sg13g2_fill_8 FILLER_0_154_224 ();
 sg13g2_fill_8 FILLER_0_154_232 ();
 sg13g2_fill_8 FILLER_0_154_240 ();
 sg13g2_fill_8 FILLER_0_154_248 ();
 sg13g2_fill_8 FILLER_0_154_256 ();
 sg13g2_fill_8 FILLER_0_154_264 ();
 sg13g2_fill_8 FILLER_0_154_272 ();
 sg13g2_fill_8 FILLER_0_154_280 ();
 sg13g2_fill_8 FILLER_0_154_288 ();
 sg13g2_fill_8 FILLER_0_154_296 ();
 sg13g2_fill_8 FILLER_0_154_304 ();
 sg13g2_fill_8 FILLER_0_154_312 ();
 sg13g2_fill_8 FILLER_0_154_320 ();
 sg13g2_fill_8 FILLER_0_154_328 ();
 sg13g2_fill_8 FILLER_0_154_336 ();
 sg13g2_fill_4 FILLER_0_154_344 ();
 sg13g2_fill_2 FILLER_0_154_353 ();
 sg13g2_fill_4 FILLER_0_154_359 ();
 sg13g2_fill_2 FILLER_0_154_363 ();
 sg13g2_fill_8 FILLER_0_154_391 ();
 sg13g2_fill_2 FILLER_0_154_399 ();
 sg13g2_fill_8 FILLER_0_154_407 ();
 sg13g2_fill_4 FILLER_0_154_415 ();
 sg13g2_fill_8 FILLER_0_154_425 ();
 sg13g2_fill_2 FILLER_0_154_433 ();
 sg13g2_fill_1 FILLER_0_154_435 ();
 sg13g2_fill_8 FILLER_0_154_439 ();
 sg13g2_fill_8 FILLER_0_154_447 ();
 sg13g2_fill_1 FILLER_0_154_455 ();
 sg13g2_fill_2 FILLER_0_154_461 ();
 sg13g2_fill_1 FILLER_0_154_463 ();
 sg13g2_fill_8 FILLER_0_154_468 ();
 sg13g2_fill_8 FILLER_0_154_476 ();
 sg13g2_fill_8 FILLER_0_154_484 ();
 sg13g2_fill_8 FILLER_0_154_492 ();
 sg13g2_fill_2 FILLER_0_154_500 ();
 sg13g2_fill_1 FILLER_0_154_502 ();
 sg13g2_fill_8 FILLER_0_154_529 ();
 sg13g2_fill_8 FILLER_0_154_537 ();
 sg13g2_fill_8 FILLER_0_154_545 ();
 sg13g2_fill_8 FILLER_0_154_553 ();
 sg13g2_fill_4 FILLER_0_154_561 ();
 sg13g2_fill_2 FILLER_0_154_565 ();
 sg13g2_fill_1 FILLER_0_154_567 ();
 sg13g2_fill_2 FILLER_0_154_573 ();
 sg13g2_fill_2 FILLER_0_154_601 ();
 sg13g2_fill_4 FILLER_0_154_629 ();
 sg13g2_fill_2 FILLER_0_154_633 ();
 sg13g2_fill_1 FILLER_0_154_635 ();
 sg13g2_fill_2 FILLER_0_154_641 ();
 sg13g2_fill_4 FILLER_0_154_647 ();
 sg13g2_fill_1 FILLER_0_154_651 ();
 sg13g2_fill_2 FILLER_0_154_657 ();
 sg13g2_fill_2 FILLER_0_154_664 ();
 sg13g2_fill_1 FILLER_0_154_666 ();
 sg13g2_fill_2 FILLER_0_154_672 ();
 sg13g2_fill_1 FILLER_0_154_674 ();
 sg13g2_fill_4 FILLER_0_154_679 ();
 sg13g2_fill_1 FILLER_0_154_683 ();
 sg13g2_fill_2 FILLER_0_154_689 ();
 sg13g2_fill_8 FILLER_0_154_696 ();
 sg13g2_fill_8 FILLER_0_154_704 ();
 sg13g2_fill_8 FILLER_0_154_712 ();
 sg13g2_fill_8 FILLER_0_154_720 ();
 sg13g2_fill_8 FILLER_0_154_728 ();
 sg13g2_fill_8 FILLER_0_154_736 ();
 sg13g2_fill_2 FILLER_0_154_749 ();
 sg13g2_fill_8 FILLER_0_154_755 ();
 sg13g2_fill_8 FILLER_0_154_763 ();
 sg13g2_fill_2 FILLER_0_154_771 ();
 sg13g2_fill_8 FILLER_0_154_777 ();
 sg13g2_fill_2 FILLER_0_154_785 ();
 sg13g2_fill_1 FILLER_0_154_787 ();
 sg13g2_fill_2 FILLER_0_154_793 ();
 sg13g2_fill_8 FILLER_0_154_821 ();
 sg13g2_fill_8 FILLER_0_154_829 ();
 sg13g2_fill_2 FILLER_0_154_837 ();
 sg13g2_fill_2 FILLER_0_154_844 ();
 sg13g2_fill_2 FILLER_0_154_851 ();
 sg13g2_fill_1 FILLER_0_154_853 ();
 sg13g2_fill_4 FILLER_0_154_858 ();
 sg13g2_fill_2 FILLER_0_154_862 ();
 sg13g2_fill_1 FILLER_0_154_864 ();
 sg13g2_fill_2 FILLER_0_154_872 ();
 sg13g2_fill_1 FILLER_0_154_874 ();
 sg13g2_fill_4 FILLER_0_154_901 ();
 sg13g2_fill_2 FILLER_0_154_905 ();
 sg13g2_fill_1 FILLER_0_154_907 ();
 sg13g2_fill_2 FILLER_0_154_929 ();
 sg13g2_fill_4 FILLER_0_154_936 ();
 sg13g2_fill_2 FILLER_0_154_940 ();
 sg13g2_fill_1 FILLER_0_154_942 ();
 sg13g2_fill_2 FILLER_0_154_947 ();
 sg13g2_fill_8 FILLER_0_154_953 ();
 sg13g2_fill_8 FILLER_0_154_966 ();
 sg13g2_fill_8 FILLER_0_154_978 ();
 sg13g2_fill_8 FILLER_0_154_986 ();
 sg13g2_fill_8 FILLER_0_154_994 ();
 sg13g2_fill_4 FILLER_0_154_1002 ();
 sg13g2_fill_4 FILLER_0_154_1011 ();
 sg13g2_fill_2 FILLER_0_154_1015 ();
 sg13g2_fill_1 FILLER_0_154_1017 ();
 sg13g2_fill_2 FILLER_0_154_1044 ();
 sg13g2_fill_8 FILLER_0_154_1052 ();
 sg13g2_fill_8 FILLER_0_154_1060 ();
 sg13g2_fill_8 FILLER_0_154_1068 ();
 sg13g2_fill_8 FILLER_0_154_1076 ();
 sg13g2_fill_1 FILLER_0_154_1084 ();
 sg13g2_fill_8 FILLER_0_154_1106 ();
 sg13g2_fill_2 FILLER_0_154_1114 ();
 sg13g2_fill_1 FILLER_0_154_1116 ();
 sg13g2_fill_2 FILLER_0_154_1122 ();
 sg13g2_fill_8 FILLER_0_154_1128 ();
 sg13g2_fill_4 FILLER_0_154_1141 ();
 sg13g2_fill_2 FILLER_0_154_1145 ();
 sg13g2_fill_4 FILLER_0_154_1153 ();
 sg13g2_fill_2 FILLER_0_154_1157 ();
 sg13g2_fill_1 FILLER_0_154_1159 ();
 sg13g2_fill_8 FILLER_0_154_1165 ();
 sg13g2_fill_8 FILLER_0_154_1173 ();
 sg13g2_fill_2 FILLER_0_154_1181 ();
 sg13g2_fill_8 FILLER_0_154_1187 ();
 sg13g2_fill_4 FILLER_0_154_1195 ();
 sg13g2_fill_2 FILLER_0_154_1199 ();
 sg13g2_fill_2 FILLER_0_154_1222 ();
 sg13g2_fill_1 FILLER_0_154_1224 ();
 sg13g2_fill_2 FILLER_0_154_1230 ();
 sg13g2_fill_1 FILLER_0_154_1232 ();
 sg13g2_fill_2 FILLER_0_154_1243 ();
 sg13g2_fill_8 FILLER_0_154_1250 ();
 sg13g2_fill_8 FILLER_0_154_1258 ();
 sg13g2_fill_8 FILLER_0_154_1266 ();
 sg13g2_fill_8 FILLER_0_154_1274 ();
 sg13g2_fill_8 FILLER_0_154_1282 ();
 sg13g2_fill_4 FILLER_0_154_1290 ();
 sg13g2_fill_2 FILLER_0_154_1294 ();
 sg13g2_fill_1 FILLER_0_154_1296 ();
 sg13g2_fill_8 FILLER_0_155_0 ();
 sg13g2_fill_8 FILLER_0_155_8 ();
 sg13g2_fill_8 FILLER_0_155_16 ();
 sg13g2_fill_8 FILLER_0_155_24 ();
 sg13g2_fill_8 FILLER_0_155_32 ();
 sg13g2_fill_8 FILLER_0_155_40 ();
 sg13g2_fill_8 FILLER_0_155_48 ();
 sg13g2_fill_8 FILLER_0_155_56 ();
 sg13g2_fill_8 FILLER_0_155_64 ();
 sg13g2_fill_8 FILLER_0_155_72 ();
 sg13g2_fill_8 FILLER_0_155_80 ();
 sg13g2_fill_8 FILLER_0_155_88 ();
 sg13g2_fill_8 FILLER_0_155_96 ();
 sg13g2_fill_8 FILLER_0_155_104 ();
 sg13g2_fill_8 FILLER_0_155_112 ();
 sg13g2_fill_8 FILLER_0_155_120 ();
 sg13g2_fill_8 FILLER_0_155_128 ();
 sg13g2_fill_8 FILLER_0_155_136 ();
 sg13g2_fill_8 FILLER_0_155_144 ();
 sg13g2_fill_8 FILLER_0_155_152 ();
 sg13g2_fill_8 FILLER_0_155_160 ();
 sg13g2_fill_8 FILLER_0_155_168 ();
 sg13g2_fill_8 FILLER_0_155_176 ();
 sg13g2_fill_8 FILLER_0_155_184 ();
 sg13g2_fill_8 FILLER_0_155_192 ();
 sg13g2_fill_8 FILLER_0_155_200 ();
 sg13g2_fill_8 FILLER_0_155_208 ();
 sg13g2_fill_8 FILLER_0_155_216 ();
 sg13g2_fill_8 FILLER_0_155_224 ();
 sg13g2_fill_8 FILLER_0_155_232 ();
 sg13g2_fill_8 FILLER_0_155_240 ();
 sg13g2_fill_8 FILLER_0_155_248 ();
 sg13g2_fill_8 FILLER_0_155_256 ();
 sg13g2_fill_8 FILLER_0_155_264 ();
 sg13g2_fill_8 FILLER_0_155_272 ();
 sg13g2_fill_8 FILLER_0_155_280 ();
 sg13g2_fill_8 FILLER_0_155_288 ();
 sg13g2_fill_8 FILLER_0_155_296 ();
 sg13g2_fill_8 FILLER_0_155_304 ();
 sg13g2_fill_8 FILLER_0_155_312 ();
 sg13g2_fill_8 FILLER_0_155_320 ();
 sg13g2_fill_4 FILLER_0_155_328 ();
 sg13g2_fill_2 FILLER_0_155_332 ();
 sg13g2_fill_1 FILLER_0_155_334 ();
 sg13g2_fill_4 FILLER_0_155_361 ();
 sg13g2_fill_2 FILLER_0_155_365 ();
 sg13g2_fill_2 FILLER_0_155_372 ();
 sg13g2_fill_8 FILLER_0_155_378 ();
 sg13g2_fill_8 FILLER_0_155_386 ();
 sg13g2_fill_8 FILLER_0_155_394 ();
 sg13g2_fill_8 FILLER_0_155_402 ();
 sg13g2_fill_2 FILLER_0_155_415 ();
 sg13g2_fill_8 FILLER_0_155_443 ();
 sg13g2_fill_2 FILLER_0_155_451 ();
 sg13g2_fill_8 FILLER_0_155_479 ();
 sg13g2_fill_8 FILLER_0_155_487 ();
 sg13g2_fill_8 FILLER_0_155_495 ();
 sg13g2_fill_2 FILLER_0_155_503 ();
 sg13g2_fill_8 FILLER_0_155_515 ();
 sg13g2_fill_4 FILLER_0_155_523 ();
 sg13g2_fill_8 FILLER_0_155_548 ();
 sg13g2_fill_4 FILLER_0_155_556 ();
 sg13g2_fill_8 FILLER_0_155_565 ();
 sg13g2_fill_8 FILLER_0_155_573 ();
 sg13g2_fill_4 FILLER_0_155_581 ();
 sg13g2_fill_2 FILLER_0_155_585 ();
 sg13g2_fill_1 FILLER_0_155_587 ();
 sg13g2_fill_8 FILLER_0_155_598 ();
 sg13g2_fill_8 FILLER_0_155_610 ();
 sg13g2_fill_8 FILLER_0_155_618 ();
 sg13g2_fill_4 FILLER_0_155_626 ();
 sg13g2_fill_1 FILLER_0_155_630 ();
 sg13g2_fill_8 FILLER_0_155_636 ();
 sg13g2_fill_8 FILLER_0_155_644 ();
 sg13g2_fill_8 FILLER_0_155_652 ();
 sg13g2_fill_8 FILLER_0_155_660 ();
 sg13g2_fill_8 FILLER_0_155_668 ();
 sg13g2_fill_2 FILLER_0_155_676 ();
 sg13g2_fill_8 FILLER_0_155_683 ();
 sg13g2_fill_8 FILLER_0_155_691 ();
 sg13g2_fill_8 FILLER_0_155_699 ();
 sg13g2_fill_8 FILLER_0_155_707 ();
 sg13g2_fill_2 FILLER_0_155_715 ();
 sg13g2_fill_4 FILLER_0_155_722 ();
 sg13g2_fill_2 FILLER_0_155_730 ();
 sg13g2_fill_8 FILLER_0_155_758 ();
 sg13g2_fill_4 FILLER_0_155_766 ();
 sg13g2_fill_8 FILLER_0_155_775 ();
 sg13g2_fill_8 FILLER_0_155_783 ();
 sg13g2_fill_4 FILLER_0_155_791 ();
 sg13g2_fill_2 FILLER_0_155_795 ();
 sg13g2_fill_1 FILLER_0_155_797 ();
 sg13g2_fill_8 FILLER_0_155_804 ();
 sg13g2_fill_8 FILLER_0_155_812 ();
 sg13g2_fill_8 FILLER_0_155_820 ();
 sg13g2_fill_4 FILLER_0_155_828 ();
 sg13g2_fill_1 FILLER_0_155_832 ();
 sg13g2_fill_8 FILLER_0_155_859 ();
 sg13g2_fill_8 FILLER_0_155_867 ();
 sg13g2_fill_8 FILLER_0_155_875 ();
 sg13g2_fill_2 FILLER_0_155_883 ();
 sg13g2_fill_1 FILLER_0_155_885 ();
 sg13g2_fill_8 FILLER_0_155_890 ();
 sg13g2_fill_4 FILLER_0_155_903 ();
 sg13g2_fill_2 FILLER_0_155_907 ();
 sg13g2_fill_2 FILLER_0_155_913 ();
 sg13g2_fill_1 FILLER_0_155_915 ();
 sg13g2_fill_2 FILLER_0_155_942 ();
 sg13g2_fill_2 FILLER_0_155_949 ();
 sg13g2_fill_1 FILLER_0_155_951 ();
 sg13g2_fill_2 FILLER_0_155_978 ();
 sg13g2_fill_4 FILLER_0_155_984 ();
 sg13g2_fill_8 FILLER_0_155_993 ();
 sg13g2_fill_8 FILLER_0_155_1001 ();
 sg13g2_fill_8 FILLER_0_155_1009 ();
 sg13g2_fill_1 FILLER_0_155_1017 ();
 sg13g2_fill_2 FILLER_0_155_1023 ();
 sg13g2_fill_2 FILLER_0_155_1030 ();
 sg13g2_fill_2 FILLER_0_155_1038 ();
 sg13g2_fill_8 FILLER_0_155_1045 ();
 sg13g2_fill_8 FILLER_0_155_1053 ();
 sg13g2_fill_4 FILLER_0_155_1061 ();
 sg13g2_fill_2 FILLER_0_155_1065 ();
 sg13g2_fill_1 FILLER_0_155_1067 ();
 sg13g2_fill_8 FILLER_0_155_1094 ();
 sg13g2_fill_4 FILLER_0_155_1107 ();
 sg13g2_fill_2 FILLER_0_155_1111 ();
 sg13g2_fill_8 FILLER_0_155_1139 ();
 sg13g2_fill_8 FILLER_0_155_1147 ();
 sg13g2_fill_8 FILLER_0_155_1155 ();
 sg13g2_fill_8 FILLER_0_155_1163 ();
 sg13g2_fill_8 FILLER_0_155_1171 ();
 sg13g2_fill_8 FILLER_0_155_1179 ();
 sg13g2_fill_8 FILLER_0_155_1187 ();
 sg13g2_fill_8 FILLER_0_155_1195 ();
 sg13g2_fill_4 FILLER_0_155_1203 ();
 sg13g2_fill_2 FILLER_0_155_1207 ();
 sg13g2_fill_8 FILLER_0_155_1235 ();
 sg13g2_fill_8 FILLER_0_155_1247 ();
 sg13g2_fill_8 FILLER_0_155_1255 ();
 sg13g2_fill_8 FILLER_0_155_1263 ();
 sg13g2_fill_8 FILLER_0_155_1271 ();
 sg13g2_fill_8 FILLER_0_155_1279 ();
 sg13g2_fill_8 FILLER_0_155_1287 ();
 sg13g2_fill_2 FILLER_0_155_1295 ();
 sg13g2_fill_8 FILLER_0_156_0 ();
 sg13g2_fill_8 FILLER_0_156_8 ();
 sg13g2_fill_8 FILLER_0_156_16 ();
 sg13g2_fill_8 FILLER_0_156_24 ();
 sg13g2_fill_8 FILLER_0_156_32 ();
 sg13g2_fill_8 FILLER_0_156_40 ();
 sg13g2_fill_8 FILLER_0_156_48 ();
 sg13g2_fill_8 FILLER_0_156_56 ();
 sg13g2_fill_8 FILLER_0_156_64 ();
 sg13g2_fill_8 FILLER_0_156_72 ();
 sg13g2_fill_8 FILLER_0_156_80 ();
 sg13g2_fill_8 FILLER_0_156_88 ();
 sg13g2_fill_8 FILLER_0_156_96 ();
 sg13g2_fill_8 FILLER_0_156_104 ();
 sg13g2_fill_8 FILLER_0_156_112 ();
 sg13g2_fill_8 FILLER_0_156_120 ();
 sg13g2_fill_8 FILLER_0_156_128 ();
 sg13g2_fill_8 FILLER_0_156_136 ();
 sg13g2_fill_8 FILLER_0_156_144 ();
 sg13g2_fill_8 FILLER_0_156_152 ();
 sg13g2_fill_8 FILLER_0_156_160 ();
 sg13g2_fill_8 FILLER_0_156_168 ();
 sg13g2_fill_8 FILLER_0_156_176 ();
 sg13g2_fill_8 FILLER_0_156_184 ();
 sg13g2_fill_8 FILLER_0_156_192 ();
 sg13g2_fill_8 FILLER_0_156_200 ();
 sg13g2_fill_8 FILLER_0_156_208 ();
 sg13g2_fill_8 FILLER_0_156_216 ();
 sg13g2_fill_8 FILLER_0_156_224 ();
 sg13g2_fill_8 FILLER_0_156_232 ();
 sg13g2_fill_8 FILLER_0_156_240 ();
 sg13g2_fill_8 FILLER_0_156_248 ();
 sg13g2_fill_8 FILLER_0_156_256 ();
 sg13g2_fill_8 FILLER_0_156_264 ();
 sg13g2_fill_8 FILLER_0_156_272 ();
 sg13g2_fill_8 FILLER_0_156_280 ();
 sg13g2_fill_8 FILLER_0_156_288 ();
 sg13g2_fill_8 FILLER_0_156_296 ();
 sg13g2_fill_8 FILLER_0_156_304 ();
 sg13g2_fill_8 FILLER_0_156_312 ();
 sg13g2_fill_8 FILLER_0_156_320 ();
 sg13g2_fill_8 FILLER_0_156_328 ();
 sg13g2_fill_8 FILLER_0_156_336 ();
 sg13g2_fill_8 FILLER_0_156_344 ();
 sg13g2_fill_8 FILLER_0_156_352 ();
 sg13g2_fill_8 FILLER_0_156_360 ();
 sg13g2_fill_8 FILLER_0_156_368 ();
 sg13g2_fill_8 FILLER_0_156_376 ();
 sg13g2_fill_8 FILLER_0_156_384 ();
 sg13g2_fill_8 FILLER_0_156_392 ();
 sg13g2_fill_4 FILLER_0_156_400 ();
 sg13g2_fill_1 FILLER_0_156_404 ();
 sg13g2_fill_2 FILLER_0_156_431 ();
 sg13g2_fill_8 FILLER_0_156_437 ();
 sg13g2_fill_8 FILLER_0_156_445 ();
 sg13g2_fill_8 FILLER_0_156_453 ();
 sg13g2_fill_8 FILLER_0_156_461 ();
 sg13g2_fill_8 FILLER_0_156_469 ();
 sg13g2_fill_4 FILLER_0_156_477 ();
 sg13g2_fill_1 FILLER_0_156_481 ();
 sg13g2_fill_8 FILLER_0_156_503 ();
 sg13g2_fill_8 FILLER_0_156_511 ();
 sg13g2_fill_4 FILLER_0_156_519 ();
 sg13g2_fill_2 FILLER_0_156_527 ();
 sg13g2_fill_2 FILLER_0_156_534 ();
 sg13g2_fill_2 FILLER_0_156_562 ();
 sg13g2_fill_2 FILLER_0_156_569 ();
 sg13g2_fill_2 FILLER_0_156_576 ();
 sg13g2_fill_8 FILLER_0_156_582 ();
 sg13g2_fill_8 FILLER_0_156_590 ();
 sg13g2_fill_8 FILLER_0_156_598 ();
 sg13g2_fill_8 FILLER_0_156_606 ();
 sg13g2_fill_8 FILLER_0_156_614 ();
 sg13g2_fill_8 FILLER_0_156_622 ();
 sg13g2_fill_8 FILLER_0_156_630 ();
 sg13g2_fill_4 FILLER_0_156_638 ();
 sg13g2_fill_2 FILLER_0_156_642 ();
 sg13g2_fill_1 FILLER_0_156_644 ();
 sg13g2_fill_2 FILLER_0_156_650 ();
 sg13g2_fill_8 FILLER_0_156_658 ();
 sg13g2_fill_8 FILLER_0_156_666 ();
 sg13g2_fill_8 FILLER_0_156_674 ();
 sg13g2_fill_8 FILLER_0_156_682 ();
 sg13g2_fill_8 FILLER_0_156_690 ();
 sg13g2_fill_2 FILLER_0_156_698 ();
 sg13g2_fill_1 FILLER_0_156_700 ();
 sg13g2_fill_8 FILLER_0_156_727 ();
 sg13g2_fill_8 FILLER_0_156_735 ();
 sg13g2_fill_8 FILLER_0_156_743 ();
 sg13g2_fill_8 FILLER_0_156_751 ();
 sg13g2_fill_4 FILLER_0_156_759 ();
 sg13g2_fill_8 FILLER_0_156_789 ();
 sg13g2_fill_8 FILLER_0_156_797 ();
 sg13g2_fill_4 FILLER_0_156_805 ();
 sg13g2_fill_1 FILLER_0_156_809 ();
 sg13g2_fill_2 FILLER_0_156_815 ();
 sg13g2_fill_4 FILLER_0_156_822 ();
 sg13g2_fill_2 FILLER_0_156_826 ();
 sg13g2_fill_1 FILLER_0_156_828 ();
 sg13g2_fill_2 FILLER_0_156_833 ();
 sg13g2_fill_1 FILLER_0_156_835 ();
 sg13g2_fill_4 FILLER_0_156_841 ();
 sg13g2_fill_2 FILLER_0_156_850 ();
 sg13g2_fill_8 FILLER_0_156_858 ();
 sg13g2_fill_8 FILLER_0_156_866 ();
 sg13g2_fill_8 FILLER_0_156_874 ();
 sg13g2_fill_8 FILLER_0_156_882 ();
 sg13g2_fill_4 FILLER_0_156_890 ();
 sg13g2_fill_4 FILLER_0_156_920 ();
 sg13g2_fill_2 FILLER_0_156_930 ();
 sg13g2_fill_2 FILLER_0_156_937 ();
 sg13g2_fill_4 FILLER_0_156_944 ();
 sg13g2_fill_2 FILLER_0_156_974 ();
 sg13g2_fill_4 FILLER_0_156_986 ();
 sg13g2_fill_2 FILLER_0_156_990 ();
 sg13g2_fill_1 FILLER_0_156_992 ();
 sg13g2_fill_4 FILLER_0_156_1019 ();
 sg13g2_fill_8 FILLER_0_156_1028 ();
 sg13g2_fill_1 FILLER_0_156_1036 ();
 sg13g2_fill_2 FILLER_0_156_1042 ();
 sg13g2_fill_8 FILLER_0_156_1048 ();
 sg13g2_fill_1 FILLER_0_156_1056 ();
 sg13g2_fill_2 FILLER_0_156_1083 ();
 sg13g2_fill_4 FILLER_0_156_1090 ();
 sg13g2_fill_2 FILLER_0_156_1094 ();
 sg13g2_fill_4 FILLER_0_156_1122 ();
 sg13g2_fill_2 FILLER_0_156_1126 ();
 sg13g2_fill_1 FILLER_0_156_1128 ();
 sg13g2_fill_8 FILLER_0_156_1135 ();
 sg13g2_fill_8 FILLER_0_156_1143 ();
 sg13g2_fill_4 FILLER_0_156_1151 ();
 sg13g2_fill_2 FILLER_0_156_1155 ();
 sg13g2_fill_2 FILLER_0_156_1162 ();
 sg13g2_fill_8 FILLER_0_156_1168 ();
 sg13g2_fill_8 FILLER_0_156_1176 ();
 sg13g2_fill_8 FILLER_0_156_1184 ();
 sg13g2_fill_2 FILLER_0_156_1192 ();
 sg13g2_fill_1 FILLER_0_156_1194 ();
 sg13g2_fill_2 FILLER_0_156_1200 ();
 sg13g2_fill_8 FILLER_0_156_1207 ();
 sg13g2_fill_8 FILLER_0_156_1215 ();
 sg13g2_fill_8 FILLER_0_156_1223 ();
 sg13g2_fill_8 FILLER_0_156_1231 ();
 sg13g2_fill_8 FILLER_0_156_1239 ();
 sg13g2_fill_8 FILLER_0_156_1247 ();
 sg13g2_fill_8 FILLER_0_156_1255 ();
 sg13g2_fill_8 FILLER_0_156_1263 ();
 sg13g2_fill_8 FILLER_0_156_1271 ();
 sg13g2_fill_8 FILLER_0_156_1279 ();
 sg13g2_fill_8 FILLER_0_156_1287 ();
 sg13g2_fill_2 FILLER_0_156_1295 ();
 sg13g2_fill_8 FILLER_0_157_0 ();
 sg13g2_fill_8 FILLER_0_157_8 ();
 sg13g2_fill_8 FILLER_0_157_16 ();
 sg13g2_fill_8 FILLER_0_157_24 ();
 sg13g2_fill_8 FILLER_0_157_32 ();
 sg13g2_fill_8 FILLER_0_157_40 ();
 sg13g2_fill_8 FILLER_0_157_48 ();
 sg13g2_fill_8 FILLER_0_157_56 ();
 sg13g2_fill_8 FILLER_0_157_64 ();
 sg13g2_fill_8 FILLER_0_157_72 ();
 sg13g2_fill_8 FILLER_0_157_80 ();
 sg13g2_fill_8 FILLER_0_157_88 ();
 sg13g2_fill_8 FILLER_0_157_96 ();
 sg13g2_fill_8 FILLER_0_157_104 ();
 sg13g2_fill_8 FILLER_0_157_112 ();
 sg13g2_fill_8 FILLER_0_157_120 ();
 sg13g2_fill_8 FILLER_0_157_128 ();
 sg13g2_fill_8 FILLER_0_157_136 ();
 sg13g2_fill_8 FILLER_0_157_144 ();
 sg13g2_fill_8 FILLER_0_157_152 ();
 sg13g2_fill_8 FILLER_0_157_160 ();
 sg13g2_fill_8 FILLER_0_157_168 ();
 sg13g2_fill_8 FILLER_0_157_176 ();
 sg13g2_fill_8 FILLER_0_157_184 ();
 sg13g2_fill_8 FILLER_0_157_192 ();
 sg13g2_fill_8 FILLER_0_157_200 ();
 sg13g2_fill_8 FILLER_0_157_208 ();
 sg13g2_fill_8 FILLER_0_157_216 ();
 sg13g2_fill_8 FILLER_0_157_224 ();
 sg13g2_fill_8 FILLER_0_157_232 ();
 sg13g2_fill_8 FILLER_0_157_240 ();
 sg13g2_fill_8 FILLER_0_157_248 ();
 sg13g2_fill_8 FILLER_0_157_256 ();
 sg13g2_fill_8 FILLER_0_157_264 ();
 sg13g2_fill_8 FILLER_0_157_272 ();
 sg13g2_fill_8 FILLER_0_157_280 ();
 sg13g2_fill_8 FILLER_0_157_288 ();
 sg13g2_fill_8 FILLER_0_157_296 ();
 sg13g2_fill_8 FILLER_0_157_304 ();
 sg13g2_fill_8 FILLER_0_157_312 ();
 sg13g2_fill_8 FILLER_0_157_320 ();
 sg13g2_fill_8 FILLER_0_157_328 ();
 sg13g2_fill_8 FILLER_0_157_336 ();
 sg13g2_fill_8 FILLER_0_157_344 ();
 sg13g2_fill_8 FILLER_0_157_352 ();
 sg13g2_fill_8 FILLER_0_157_360 ();
 sg13g2_fill_8 FILLER_0_157_368 ();
 sg13g2_fill_8 FILLER_0_157_376 ();
 sg13g2_fill_8 FILLER_0_157_384 ();
 sg13g2_fill_8 FILLER_0_157_392 ();
 sg13g2_fill_4 FILLER_0_157_400 ();
 sg13g2_fill_2 FILLER_0_157_404 ();
 sg13g2_fill_1 FILLER_0_157_406 ();
 sg13g2_fill_2 FILLER_0_157_412 ();
 sg13g2_fill_2 FILLER_0_157_418 ();
 sg13g2_fill_1 FILLER_0_157_420 ();
 sg13g2_fill_8 FILLER_0_157_426 ();
 sg13g2_fill_8 FILLER_0_157_434 ();
 sg13g2_fill_4 FILLER_0_157_442 ();
 sg13g2_fill_2 FILLER_0_157_446 ();
 sg13g2_fill_1 FILLER_0_157_448 ();
 sg13g2_fill_2 FILLER_0_157_454 ();
 sg13g2_fill_2 FILLER_0_157_482 ();
 sg13g2_fill_4 FILLER_0_157_505 ();
 sg13g2_fill_1 FILLER_0_157_509 ();
 sg13g2_fill_8 FILLER_0_157_536 ();
 sg13g2_fill_8 FILLER_0_157_549 ();
 sg13g2_fill_8 FILLER_0_157_557 ();
 sg13g2_fill_8 FILLER_0_157_565 ();
 sg13g2_fill_8 FILLER_0_157_573 ();
 sg13g2_fill_8 FILLER_0_157_581 ();
 sg13g2_fill_8 FILLER_0_157_610 ();
 sg13g2_fill_1 FILLER_0_157_618 ();
 sg13g2_fill_8 FILLER_0_157_624 ();
 sg13g2_fill_1 FILLER_0_157_632 ();
 sg13g2_fill_4 FILLER_0_157_638 ();
 sg13g2_fill_4 FILLER_0_157_647 ();
 sg13g2_fill_2 FILLER_0_157_651 ();
 sg13g2_fill_8 FILLER_0_157_657 ();
 sg13g2_fill_1 FILLER_0_157_665 ();
 sg13g2_fill_8 FILLER_0_157_671 ();
 sg13g2_fill_1 FILLER_0_157_679 ();
 sg13g2_fill_4 FILLER_0_157_706 ();
 sg13g2_fill_2 FILLER_0_157_710 ();
 sg13g2_fill_1 FILLER_0_157_712 ();
 sg13g2_fill_2 FILLER_0_157_734 ();
 sg13g2_fill_8 FILLER_0_157_741 ();
 sg13g2_fill_8 FILLER_0_157_749 ();
 sg13g2_fill_8 FILLER_0_157_757 ();
 sg13g2_fill_2 FILLER_0_157_769 ();
 sg13g2_fill_8 FILLER_0_157_775 ();
 sg13g2_fill_4 FILLER_0_157_783 ();
 sg13g2_fill_8 FILLER_0_157_792 ();
 sg13g2_fill_8 FILLER_0_157_800 ();
 sg13g2_fill_4 FILLER_0_157_808 ();
 sg13g2_fill_1 FILLER_0_157_812 ();
 sg13g2_fill_2 FILLER_0_157_839 ();
 sg13g2_fill_8 FILLER_0_157_862 ();
 sg13g2_fill_8 FILLER_0_157_870 ();
 sg13g2_fill_8 FILLER_0_157_878 ();
 sg13g2_fill_8 FILLER_0_157_886 ();
 sg13g2_fill_8 FILLER_0_157_894 ();
 sg13g2_fill_8 FILLER_0_157_902 ();
 sg13g2_fill_4 FILLER_0_157_910 ();
 sg13g2_fill_1 FILLER_0_157_914 ();
 sg13g2_fill_2 FILLER_0_157_919 ();
 sg13g2_fill_8 FILLER_0_157_926 ();
 sg13g2_fill_8 FILLER_0_157_934 ();
 sg13g2_fill_8 FILLER_0_157_942 ();
 sg13g2_fill_1 FILLER_0_157_950 ();
 sg13g2_fill_4 FILLER_0_157_956 ();
 sg13g2_fill_2 FILLER_0_157_960 ();
 sg13g2_fill_1 FILLER_0_157_962 ();
 sg13g2_fill_2 FILLER_0_157_984 ();
 sg13g2_fill_8 FILLER_0_157_991 ();
 sg13g2_fill_8 FILLER_0_157_999 ();
 sg13g2_fill_8 FILLER_0_157_1007 ();
 sg13g2_fill_1 FILLER_0_157_1015 ();
 sg13g2_fill_2 FILLER_0_157_1021 ();
 sg13g2_fill_8 FILLER_0_157_1027 ();
 sg13g2_fill_8 FILLER_0_157_1035 ();
 sg13g2_fill_8 FILLER_0_157_1043 ();
 sg13g2_fill_4 FILLER_0_157_1051 ();
 sg13g2_fill_2 FILLER_0_157_1055 ();
 sg13g2_fill_1 FILLER_0_157_1057 ();
 sg13g2_fill_2 FILLER_0_157_1065 ();
 sg13g2_fill_2 FILLER_0_157_1072 ();
 sg13g2_fill_2 FILLER_0_157_1078 ();
 sg13g2_fill_1 FILLER_0_157_1080 ();
 sg13g2_fill_2 FILLER_0_157_1087 ();
 sg13g2_fill_8 FILLER_0_157_1094 ();
 sg13g2_fill_1 FILLER_0_157_1102 ();
 sg13g2_fill_8 FILLER_0_157_1107 ();
 sg13g2_fill_4 FILLER_0_157_1115 ();
 sg13g2_fill_2 FILLER_0_157_1124 ();
 sg13g2_fill_8 FILLER_0_157_1134 ();
 sg13g2_fill_8 FILLER_0_157_1142 ();
 sg13g2_fill_2 FILLER_0_157_1150 ();
 sg13g2_fill_1 FILLER_0_157_1152 ();
 sg13g2_fill_4 FILLER_0_157_1179 ();
 sg13g2_fill_2 FILLER_0_157_1187 ();
 sg13g2_fill_8 FILLER_0_157_1194 ();
 sg13g2_fill_8 FILLER_0_157_1202 ();
 sg13g2_fill_8 FILLER_0_157_1210 ();
 sg13g2_fill_8 FILLER_0_157_1218 ();
 sg13g2_fill_8 FILLER_0_157_1226 ();
 sg13g2_fill_8 FILLER_0_157_1234 ();
 sg13g2_fill_8 FILLER_0_157_1242 ();
 sg13g2_fill_8 FILLER_0_157_1250 ();
 sg13g2_fill_8 FILLER_0_157_1258 ();
 sg13g2_fill_8 FILLER_0_157_1266 ();
 sg13g2_fill_8 FILLER_0_157_1274 ();
 sg13g2_fill_8 FILLER_0_157_1282 ();
 sg13g2_fill_4 FILLER_0_157_1290 ();
 sg13g2_fill_2 FILLER_0_157_1294 ();
 sg13g2_fill_1 FILLER_0_157_1296 ();
 sg13g2_fill_8 FILLER_0_158_0 ();
 sg13g2_fill_8 FILLER_0_158_8 ();
 sg13g2_fill_8 FILLER_0_158_16 ();
 sg13g2_fill_8 FILLER_0_158_24 ();
 sg13g2_fill_8 FILLER_0_158_32 ();
 sg13g2_fill_8 FILLER_0_158_40 ();
 sg13g2_fill_8 FILLER_0_158_48 ();
 sg13g2_fill_8 FILLER_0_158_56 ();
 sg13g2_fill_8 FILLER_0_158_64 ();
 sg13g2_fill_8 FILLER_0_158_72 ();
 sg13g2_fill_8 FILLER_0_158_80 ();
 sg13g2_fill_8 FILLER_0_158_88 ();
 sg13g2_fill_8 FILLER_0_158_96 ();
 sg13g2_fill_8 FILLER_0_158_104 ();
 sg13g2_fill_8 FILLER_0_158_112 ();
 sg13g2_fill_8 FILLER_0_158_120 ();
 sg13g2_fill_8 FILLER_0_158_128 ();
 sg13g2_fill_8 FILLER_0_158_136 ();
 sg13g2_fill_8 FILLER_0_158_144 ();
 sg13g2_fill_8 FILLER_0_158_152 ();
 sg13g2_fill_8 FILLER_0_158_160 ();
 sg13g2_fill_8 FILLER_0_158_168 ();
 sg13g2_fill_8 FILLER_0_158_176 ();
 sg13g2_fill_8 FILLER_0_158_184 ();
 sg13g2_fill_8 FILLER_0_158_192 ();
 sg13g2_fill_8 FILLER_0_158_200 ();
 sg13g2_fill_8 FILLER_0_158_208 ();
 sg13g2_fill_8 FILLER_0_158_216 ();
 sg13g2_fill_8 FILLER_0_158_224 ();
 sg13g2_fill_8 FILLER_0_158_232 ();
 sg13g2_fill_8 FILLER_0_158_240 ();
 sg13g2_fill_8 FILLER_0_158_248 ();
 sg13g2_fill_8 FILLER_0_158_256 ();
 sg13g2_fill_8 FILLER_0_158_264 ();
 sg13g2_fill_8 FILLER_0_158_272 ();
 sg13g2_fill_8 FILLER_0_158_280 ();
 sg13g2_fill_8 FILLER_0_158_288 ();
 sg13g2_fill_8 FILLER_0_158_296 ();
 sg13g2_fill_8 FILLER_0_158_304 ();
 sg13g2_fill_8 FILLER_0_158_312 ();
 sg13g2_fill_8 FILLER_0_158_320 ();
 sg13g2_fill_8 FILLER_0_158_328 ();
 sg13g2_fill_8 FILLER_0_158_336 ();
 sg13g2_fill_8 FILLER_0_158_344 ();
 sg13g2_fill_8 FILLER_0_158_352 ();
 sg13g2_fill_8 FILLER_0_158_360 ();
 sg13g2_fill_8 FILLER_0_158_368 ();
 sg13g2_fill_8 FILLER_0_158_376 ();
 sg13g2_fill_8 FILLER_0_158_384 ();
 sg13g2_fill_8 FILLER_0_158_392 ();
 sg13g2_fill_8 FILLER_0_158_400 ();
 sg13g2_fill_8 FILLER_0_158_408 ();
 sg13g2_fill_8 FILLER_0_158_416 ();
 sg13g2_fill_8 FILLER_0_158_424 ();
 sg13g2_fill_8 FILLER_0_158_432 ();
 sg13g2_fill_8 FILLER_0_158_440 ();
 sg13g2_fill_8 FILLER_0_158_448 ();
 sg13g2_fill_1 FILLER_0_158_456 ();
 sg13g2_fill_2 FILLER_0_158_483 ();
 sg13g2_fill_4 FILLER_0_158_511 ();
 sg13g2_fill_2 FILLER_0_158_515 ();
 sg13g2_fill_2 FILLER_0_158_522 ();
 sg13g2_fill_1 FILLER_0_158_524 ();
 sg13g2_fill_8 FILLER_0_158_529 ();
 sg13g2_fill_4 FILLER_0_158_537 ();
 sg13g2_fill_2 FILLER_0_158_541 ();
 sg13g2_fill_1 FILLER_0_158_543 ();
 sg13g2_fill_2 FILLER_0_158_570 ();
 sg13g2_fill_1 FILLER_0_158_572 ();
 sg13g2_fill_2 FILLER_0_158_599 ();
 sg13g2_fill_8 FILLER_0_158_606 ();
 sg13g2_fill_8 FILLER_0_158_614 ();
 sg13g2_fill_8 FILLER_0_158_622 ();
 sg13g2_fill_1 FILLER_0_158_630 ();
 sg13g2_fill_2 FILLER_0_158_636 ();
 sg13g2_fill_2 FILLER_0_158_642 ();
 sg13g2_fill_2 FILLER_0_158_670 ();
 sg13g2_fill_2 FILLER_0_158_680 ();
 sg13g2_fill_2 FILLER_0_158_687 ();
 sg13g2_fill_4 FILLER_0_158_693 ();
 sg13g2_fill_4 FILLER_0_158_705 ();
 sg13g2_fill_8 FILLER_0_158_714 ();
 sg13g2_fill_4 FILLER_0_158_722 ();
 sg13g2_fill_2 FILLER_0_158_726 ();
 sg13g2_fill_1 FILLER_0_158_728 ();
 sg13g2_fill_4 FILLER_0_158_735 ();
 sg13g2_fill_8 FILLER_0_158_744 ();
 sg13g2_fill_8 FILLER_0_158_752 ();
 sg13g2_fill_2 FILLER_0_158_760 ();
 sg13g2_fill_8 FILLER_0_158_767 ();
 sg13g2_fill_4 FILLER_0_158_775 ();
 sg13g2_fill_1 FILLER_0_158_779 ();
 sg13g2_fill_8 FILLER_0_158_785 ();
 sg13g2_fill_8 FILLER_0_158_793 ();
 sg13g2_fill_8 FILLER_0_158_801 ();
 sg13g2_fill_8 FILLER_0_158_809 ();
 sg13g2_fill_2 FILLER_0_158_817 ();
 sg13g2_fill_1 FILLER_0_158_819 ();
 sg13g2_fill_8 FILLER_0_158_825 ();
 sg13g2_fill_8 FILLER_0_158_833 ();
 sg13g2_fill_8 FILLER_0_158_841 ();
 sg13g2_fill_8 FILLER_0_158_849 ();
 sg13g2_fill_2 FILLER_0_158_857 ();
 sg13g2_fill_2 FILLER_0_158_867 ();
 sg13g2_fill_4 FILLER_0_158_874 ();
 sg13g2_fill_2 FILLER_0_158_878 ();
 sg13g2_fill_2 FILLER_0_158_884 ();
 sg13g2_fill_8 FILLER_0_158_890 ();
 sg13g2_fill_8 FILLER_0_158_898 ();
 sg13g2_fill_1 FILLER_0_158_906 ();
 sg13g2_fill_8 FILLER_0_158_912 ();
 sg13g2_fill_8 FILLER_0_158_920 ();
 sg13g2_fill_8 FILLER_0_158_928 ();
 sg13g2_fill_8 FILLER_0_158_936 ();
 sg13g2_fill_8 FILLER_0_158_944 ();
 sg13g2_fill_2 FILLER_0_158_952 ();
 sg13g2_fill_2 FILLER_0_158_959 ();
 sg13g2_fill_1 FILLER_0_158_961 ();
 sg13g2_fill_2 FILLER_0_158_966 ();
 sg13g2_fill_8 FILLER_0_158_972 ();
 sg13g2_fill_8 FILLER_0_158_980 ();
 sg13g2_fill_8 FILLER_0_158_988 ();
 sg13g2_fill_8 FILLER_0_158_996 ();
 sg13g2_fill_8 FILLER_0_158_1004 ();
 sg13g2_fill_8 FILLER_0_158_1038 ();
 sg13g2_fill_8 FILLER_0_158_1046 ();
 sg13g2_fill_4 FILLER_0_158_1054 ();
 sg13g2_fill_2 FILLER_0_158_1058 ();
 sg13g2_fill_2 FILLER_0_158_1065 ();
 sg13g2_fill_2 FILLER_0_158_1072 ();
 sg13g2_fill_8 FILLER_0_158_1079 ();
 sg13g2_fill_8 FILLER_0_158_1087 ();
 sg13g2_fill_8 FILLER_0_158_1095 ();
 sg13g2_fill_8 FILLER_0_158_1103 ();
 sg13g2_fill_8 FILLER_0_158_1111 ();
 sg13g2_fill_8 FILLER_0_158_1119 ();
 sg13g2_fill_4 FILLER_0_158_1127 ();
 sg13g2_fill_1 FILLER_0_158_1131 ();
 sg13g2_fill_2 FILLER_0_158_1137 ();
 sg13g2_fill_8 FILLER_0_158_1144 ();
 sg13g2_fill_4 FILLER_0_158_1152 ();
 sg13g2_fill_1 FILLER_0_158_1156 ();
 sg13g2_fill_4 FILLER_0_158_1167 ();
 sg13g2_fill_1 FILLER_0_158_1171 ();
 sg13g2_fill_2 FILLER_0_158_1178 ();
 sg13g2_fill_8 FILLER_0_158_1185 ();
 sg13g2_fill_8 FILLER_0_158_1193 ();
 sg13g2_fill_2 FILLER_0_158_1201 ();
 sg13g2_fill_1 FILLER_0_158_1203 ();
 sg13g2_fill_4 FILLER_0_158_1230 ();
 sg13g2_fill_1 FILLER_0_158_1234 ();
 sg13g2_fill_8 FILLER_0_158_1245 ();
 sg13g2_fill_8 FILLER_0_158_1253 ();
 sg13g2_fill_8 FILLER_0_158_1261 ();
 sg13g2_fill_8 FILLER_0_158_1269 ();
 sg13g2_fill_8 FILLER_0_158_1277 ();
 sg13g2_fill_8 FILLER_0_158_1285 ();
 sg13g2_fill_4 FILLER_0_158_1293 ();
 sg13g2_fill_8 FILLER_0_159_0 ();
 sg13g2_fill_8 FILLER_0_159_8 ();
 sg13g2_fill_8 FILLER_0_159_16 ();
 sg13g2_fill_8 FILLER_0_159_24 ();
 sg13g2_fill_8 FILLER_0_159_32 ();
 sg13g2_fill_8 FILLER_0_159_40 ();
 sg13g2_fill_8 FILLER_0_159_48 ();
 sg13g2_fill_8 FILLER_0_159_56 ();
 sg13g2_fill_8 FILLER_0_159_64 ();
 sg13g2_fill_8 FILLER_0_159_72 ();
 sg13g2_fill_8 FILLER_0_159_80 ();
 sg13g2_fill_8 FILLER_0_159_88 ();
 sg13g2_fill_8 FILLER_0_159_96 ();
 sg13g2_fill_8 FILLER_0_159_104 ();
 sg13g2_fill_8 FILLER_0_159_112 ();
 sg13g2_fill_8 FILLER_0_159_120 ();
 sg13g2_fill_8 FILLER_0_159_128 ();
 sg13g2_fill_8 FILLER_0_159_136 ();
 sg13g2_fill_8 FILLER_0_159_144 ();
 sg13g2_fill_8 FILLER_0_159_152 ();
 sg13g2_fill_8 FILLER_0_159_160 ();
 sg13g2_fill_8 FILLER_0_159_168 ();
 sg13g2_fill_8 FILLER_0_159_176 ();
 sg13g2_fill_8 FILLER_0_159_184 ();
 sg13g2_fill_8 FILLER_0_159_192 ();
 sg13g2_fill_8 FILLER_0_159_200 ();
 sg13g2_fill_8 FILLER_0_159_208 ();
 sg13g2_fill_8 FILLER_0_159_216 ();
 sg13g2_fill_8 FILLER_0_159_224 ();
 sg13g2_fill_8 FILLER_0_159_232 ();
 sg13g2_fill_8 FILLER_0_159_240 ();
 sg13g2_fill_8 FILLER_0_159_248 ();
 sg13g2_fill_8 FILLER_0_159_256 ();
 sg13g2_fill_8 FILLER_0_159_264 ();
 sg13g2_fill_8 FILLER_0_159_272 ();
 sg13g2_fill_8 FILLER_0_159_280 ();
 sg13g2_fill_8 FILLER_0_159_288 ();
 sg13g2_fill_8 FILLER_0_159_296 ();
 sg13g2_fill_8 FILLER_0_159_304 ();
 sg13g2_fill_8 FILLER_0_159_312 ();
 sg13g2_fill_8 FILLER_0_159_320 ();
 sg13g2_fill_8 FILLER_0_159_328 ();
 sg13g2_fill_8 FILLER_0_159_336 ();
 sg13g2_fill_8 FILLER_0_159_344 ();
 sg13g2_fill_8 FILLER_0_159_352 ();
 sg13g2_fill_8 FILLER_0_159_360 ();
 sg13g2_fill_8 FILLER_0_159_368 ();
 sg13g2_fill_8 FILLER_0_159_376 ();
 sg13g2_fill_8 FILLER_0_159_384 ();
 sg13g2_fill_8 FILLER_0_159_392 ();
 sg13g2_fill_8 FILLER_0_159_400 ();
 sg13g2_fill_8 FILLER_0_159_408 ();
 sg13g2_fill_8 FILLER_0_159_416 ();
 sg13g2_fill_8 FILLER_0_159_424 ();
 sg13g2_fill_8 FILLER_0_159_432 ();
 sg13g2_fill_8 FILLER_0_159_440 ();
 sg13g2_fill_8 FILLER_0_159_448 ();
 sg13g2_fill_1 FILLER_0_159_456 ();
 sg13g2_fill_2 FILLER_0_159_462 ();
 sg13g2_fill_2 FILLER_0_159_468 ();
 sg13g2_fill_4 FILLER_0_159_474 ();
 sg13g2_fill_1 FILLER_0_159_478 ();
 sg13g2_fill_4 FILLER_0_159_484 ();
 sg13g2_fill_1 FILLER_0_159_488 ();
 sg13g2_fill_8 FILLER_0_159_493 ();
 sg13g2_fill_8 FILLER_0_159_501 ();
 sg13g2_fill_2 FILLER_0_159_509 ();
 sg13g2_fill_8 FILLER_0_159_519 ();
 sg13g2_fill_8 FILLER_0_159_527 ();
 sg13g2_fill_8 FILLER_0_159_535 ();
 sg13g2_fill_4 FILLER_0_159_543 ();
 sg13g2_fill_8 FILLER_0_159_551 ();
 sg13g2_fill_8 FILLER_0_159_559 ();
 sg13g2_fill_2 FILLER_0_159_567 ();
 sg13g2_fill_1 FILLER_0_159_569 ();
 sg13g2_fill_8 FILLER_0_159_596 ();
 sg13g2_fill_1 FILLER_0_159_604 ();
 sg13g2_fill_8 FILLER_0_159_610 ();
 sg13g2_fill_4 FILLER_0_159_618 ();
 sg13g2_fill_8 FILLER_0_159_648 ();
 sg13g2_fill_1 FILLER_0_159_656 ();
 sg13g2_fill_8 FILLER_0_159_678 ();
 sg13g2_fill_8 FILLER_0_159_686 ();
 sg13g2_fill_8 FILLER_0_159_694 ();
 sg13g2_fill_4 FILLER_0_159_707 ();
 sg13g2_fill_2 FILLER_0_159_711 ();
 sg13g2_fill_4 FILLER_0_159_717 ();
 sg13g2_fill_8 FILLER_0_159_726 ();
 sg13g2_fill_4 FILLER_0_159_734 ();
 sg13g2_fill_2 FILLER_0_159_738 ();
 sg13g2_fill_2 FILLER_0_159_748 ();
 sg13g2_fill_1 FILLER_0_159_750 ();
 sg13g2_fill_2 FILLER_0_159_757 ();
 sg13g2_fill_1 FILLER_0_159_759 ();
 sg13g2_fill_2 FILLER_0_159_765 ();
 sg13g2_fill_1 FILLER_0_159_767 ();
 sg13g2_fill_4 FILLER_0_159_774 ();
 sg13g2_fill_2 FILLER_0_159_782 ();
 sg13g2_fill_1 FILLER_0_159_784 ();
 sg13g2_fill_2 FILLER_0_159_811 ();
 sg13g2_fill_4 FILLER_0_159_818 ();
 sg13g2_fill_1 FILLER_0_159_822 ();
 sg13g2_fill_8 FILLER_0_159_828 ();
 sg13g2_fill_1 FILLER_0_159_836 ();
 sg13g2_fill_4 FILLER_0_159_845 ();
 sg13g2_fill_1 FILLER_0_159_849 ();
 sg13g2_fill_4 FILLER_0_159_856 ();
 sg13g2_fill_2 FILLER_0_159_866 ();
 sg13g2_fill_2 FILLER_0_159_894 ();
 sg13g2_fill_8 FILLER_0_159_902 ();
 sg13g2_fill_8 FILLER_0_159_910 ();
 sg13g2_fill_4 FILLER_0_159_918 ();
 sg13g2_fill_8 FILLER_0_159_927 ();
 sg13g2_fill_8 FILLER_0_159_935 ();
 sg13g2_fill_8 FILLER_0_159_943 ();
 sg13g2_fill_8 FILLER_0_159_951 ();
 sg13g2_fill_4 FILLER_0_159_959 ();
 sg13g2_fill_2 FILLER_0_159_968 ();
 sg13g2_fill_2 FILLER_0_159_996 ();
 sg13g2_fill_4 FILLER_0_159_1003 ();
 sg13g2_fill_2 FILLER_0_159_1007 ();
 sg13g2_fill_1 FILLER_0_159_1009 ();
 sg13g2_fill_8 FILLER_0_159_1015 ();
 sg13g2_fill_2 FILLER_0_159_1023 ();
 sg13g2_fill_2 FILLER_0_159_1030 ();
 sg13g2_fill_8 FILLER_0_159_1038 ();
 sg13g2_fill_8 FILLER_0_159_1046 ();
 sg13g2_fill_1 FILLER_0_159_1054 ();
 sg13g2_fill_2 FILLER_0_159_1060 ();
 sg13g2_fill_2 FILLER_0_159_1066 ();
 sg13g2_fill_2 FILLER_0_159_1073 ();
 sg13g2_fill_1 FILLER_0_159_1075 ();
 sg13g2_fill_2 FILLER_0_159_1082 ();
 sg13g2_fill_8 FILLER_0_159_1089 ();
 sg13g2_fill_4 FILLER_0_159_1097 ();
 sg13g2_fill_2 FILLER_0_159_1101 ();
 sg13g2_fill_8 FILLER_0_159_1107 ();
 sg13g2_fill_8 FILLER_0_159_1115 ();
 sg13g2_fill_2 FILLER_0_159_1123 ();
 sg13g2_fill_2 FILLER_0_159_1131 ();
 sg13g2_fill_8 FILLER_0_159_1139 ();
 sg13g2_fill_4 FILLER_0_159_1147 ();
 sg13g2_fill_2 FILLER_0_159_1156 ();
 sg13g2_fill_8 FILLER_0_159_1162 ();
 sg13g2_fill_8 FILLER_0_159_1170 ();
 sg13g2_fill_2 FILLER_0_159_1182 ();
 sg13g2_fill_2 FILLER_0_159_1189 ();
 sg13g2_fill_2 FILLER_0_159_1217 ();
 sg13g2_fill_1 FILLER_0_159_1219 ();
 sg13g2_fill_2 FILLER_0_159_1225 ();
 sg13g2_fill_8 FILLER_0_159_1253 ();
 sg13g2_fill_8 FILLER_0_159_1261 ();
 sg13g2_fill_8 FILLER_0_159_1269 ();
 sg13g2_fill_8 FILLER_0_159_1277 ();
 sg13g2_fill_8 FILLER_0_159_1285 ();
 sg13g2_fill_4 FILLER_0_159_1293 ();
 sg13g2_fill_8 FILLER_0_160_0 ();
 sg13g2_fill_8 FILLER_0_160_8 ();
 sg13g2_fill_8 FILLER_0_160_16 ();
 sg13g2_fill_8 FILLER_0_160_24 ();
 sg13g2_fill_8 FILLER_0_160_32 ();
 sg13g2_fill_8 FILLER_0_160_40 ();
 sg13g2_fill_8 FILLER_0_160_48 ();
 sg13g2_fill_8 FILLER_0_160_56 ();
 sg13g2_fill_8 FILLER_0_160_64 ();
 sg13g2_fill_8 FILLER_0_160_72 ();
 sg13g2_fill_8 FILLER_0_160_80 ();
 sg13g2_fill_8 FILLER_0_160_88 ();
 sg13g2_fill_8 FILLER_0_160_96 ();
 sg13g2_fill_8 FILLER_0_160_104 ();
 sg13g2_fill_8 FILLER_0_160_112 ();
 sg13g2_fill_8 FILLER_0_160_120 ();
 sg13g2_fill_8 FILLER_0_160_128 ();
 sg13g2_fill_8 FILLER_0_160_136 ();
 sg13g2_fill_8 FILLER_0_160_144 ();
 sg13g2_fill_8 FILLER_0_160_152 ();
 sg13g2_fill_8 FILLER_0_160_160 ();
 sg13g2_fill_8 FILLER_0_160_168 ();
 sg13g2_fill_8 FILLER_0_160_176 ();
 sg13g2_fill_8 FILLER_0_160_184 ();
 sg13g2_fill_8 FILLER_0_160_192 ();
 sg13g2_fill_8 FILLER_0_160_200 ();
 sg13g2_fill_8 FILLER_0_160_208 ();
 sg13g2_fill_8 FILLER_0_160_216 ();
 sg13g2_fill_8 FILLER_0_160_224 ();
 sg13g2_fill_8 FILLER_0_160_232 ();
 sg13g2_fill_8 FILLER_0_160_240 ();
 sg13g2_fill_8 FILLER_0_160_248 ();
 sg13g2_fill_8 FILLER_0_160_256 ();
 sg13g2_fill_8 FILLER_0_160_264 ();
 sg13g2_fill_8 FILLER_0_160_272 ();
 sg13g2_fill_8 FILLER_0_160_280 ();
 sg13g2_fill_8 FILLER_0_160_288 ();
 sg13g2_fill_8 FILLER_0_160_296 ();
 sg13g2_fill_8 FILLER_0_160_304 ();
 sg13g2_fill_8 FILLER_0_160_312 ();
 sg13g2_fill_8 FILLER_0_160_320 ();
 sg13g2_fill_8 FILLER_0_160_328 ();
 sg13g2_fill_8 FILLER_0_160_336 ();
 sg13g2_fill_8 FILLER_0_160_344 ();
 sg13g2_fill_8 FILLER_0_160_352 ();
 sg13g2_fill_8 FILLER_0_160_360 ();
 sg13g2_fill_8 FILLER_0_160_368 ();
 sg13g2_fill_8 FILLER_0_160_376 ();
 sg13g2_fill_8 FILLER_0_160_384 ();
 sg13g2_fill_8 FILLER_0_160_392 ();
 sg13g2_fill_8 FILLER_0_160_400 ();
 sg13g2_fill_8 FILLER_0_160_408 ();
 sg13g2_fill_8 FILLER_0_160_416 ();
 sg13g2_fill_8 FILLER_0_160_424 ();
 sg13g2_fill_8 FILLER_0_160_432 ();
 sg13g2_fill_8 FILLER_0_160_440 ();
 sg13g2_fill_8 FILLER_0_160_448 ();
 sg13g2_fill_8 FILLER_0_160_456 ();
 sg13g2_fill_8 FILLER_0_160_464 ();
 sg13g2_fill_8 FILLER_0_160_472 ();
 sg13g2_fill_8 FILLER_0_160_480 ();
 sg13g2_fill_8 FILLER_0_160_488 ();
 sg13g2_fill_8 FILLER_0_160_496 ();
 sg13g2_fill_8 FILLER_0_160_504 ();
 sg13g2_fill_8 FILLER_0_160_512 ();
 sg13g2_fill_8 FILLER_0_160_520 ();
 sg13g2_fill_8 FILLER_0_160_528 ();
 sg13g2_fill_8 FILLER_0_160_536 ();
 sg13g2_fill_8 FILLER_0_160_544 ();
 sg13g2_fill_8 FILLER_0_160_552 ();
 sg13g2_fill_8 FILLER_0_160_560 ();
 sg13g2_fill_4 FILLER_0_160_568 ();
 sg13g2_fill_1 FILLER_0_160_572 ();
 sg13g2_fill_2 FILLER_0_160_578 ();
 sg13g2_fill_8 FILLER_0_160_584 ();
 sg13g2_fill_8 FILLER_0_160_592 ();
 sg13g2_fill_8 FILLER_0_160_600 ();
 sg13g2_fill_8 FILLER_0_160_608 ();
 sg13g2_fill_8 FILLER_0_160_616 ();
 sg13g2_fill_8 FILLER_0_160_624 ();
 sg13g2_fill_8 FILLER_0_160_632 ();
 sg13g2_fill_4 FILLER_0_160_640 ();
 sg13g2_fill_1 FILLER_0_160_644 ();
 sg13g2_fill_2 FILLER_0_160_649 ();
 sg13g2_fill_8 FILLER_0_160_661 ();
 sg13g2_fill_8 FILLER_0_160_669 ();
 sg13g2_fill_8 FILLER_0_160_677 ();
 sg13g2_fill_8 FILLER_0_160_685 ();
 sg13g2_fill_2 FILLER_0_160_693 ();
 sg13g2_fill_2 FILLER_0_160_700 ();
 sg13g2_fill_2 FILLER_0_160_728 ();
 sg13g2_fill_8 FILLER_0_160_740 ();
 sg13g2_fill_2 FILLER_0_160_748 ();
 sg13g2_fill_1 FILLER_0_160_750 ();
 sg13g2_fill_2 FILLER_0_160_777 ();
 sg13g2_fill_8 FILLER_0_160_785 ();
 sg13g2_fill_4 FILLER_0_160_793 ();
 sg13g2_fill_2 FILLER_0_160_797 ();
 sg13g2_fill_2 FILLER_0_160_806 ();
 sg13g2_fill_4 FILLER_0_160_813 ();
 sg13g2_fill_2 FILLER_0_160_817 ();
 sg13g2_fill_2 FILLER_0_160_824 ();
 sg13g2_fill_2 FILLER_0_160_852 ();
 sg13g2_fill_4 FILLER_0_160_858 ();
 sg13g2_fill_2 FILLER_0_160_867 ();
 sg13g2_fill_2 FILLER_0_160_874 ();
 sg13g2_fill_1 FILLER_0_160_876 ();
 sg13g2_fill_4 FILLER_0_160_882 ();
 sg13g2_fill_1 FILLER_0_160_886 ();
 sg13g2_fill_4 FILLER_0_160_892 ();
 sg13g2_fill_2 FILLER_0_160_896 ();
 sg13g2_fill_4 FILLER_0_160_904 ();
 sg13g2_fill_2 FILLER_0_160_908 ();
 sg13g2_fill_1 FILLER_0_160_910 ();
 sg13g2_fill_8 FILLER_0_160_937 ();
 sg13g2_fill_8 FILLER_0_160_945 ();
 sg13g2_fill_4 FILLER_0_160_953 ();
 sg13g2_fill_2 FILLER_0_160_957 ();
 sg13g2_fill_1 FILLER_0_160_959 ();
 sg13g2_fill_2 FILLER_0_160_986 ();
 sg13g2_fill_2 FILLER_0_160_993 ();
 sg13g2_fill_4 FILLER_0_160_1000 ();
 sg13g2_fill_2 FILLER_0_160_1004 ();
 sg13g2_fill_8 FILLER_0_160_1010 ();
 sg13g2_fill_8 FILLER_0_160_1022 ();
 sg13g2_fill_8 FILLER_0_160_1030 ();
 sg13g2_fill_4 FILLER_0_160_1038 ();
 sg13g2_fill_2 FILLER_0_160_1042 ();
 sg13g2_fill_8 FILLER_0_160_1049 ();
 sg13g2_fill_8 FILLER_0_160_1057 ();
 sg13g2_fill_2 FILLER_0_160_1065 ();
 sg13g2_fill_8 FILLER_0_160_1072 ();
 sg13g2_fill_2 FILLER_0_160_1080 ();
 sg13g2_fill_8 FILLER_0_160_1087 ();
 sg13g2_fill_4 FILLER_0_160_1095 ();
 sg13g2_fill_2 FILLER_0_160_1104 ();
 sg13g2_fill_2 FILLER_0_160_1132 ();
 sg13g2_fill_4 FILLER_0_160_1140 ();
 sg13g2_fill_2 FILLER_0_160_1144 ();
 sg13g2_fill_1 FILLER_0_160_1146 ();
 sg13g2_fill_2 FILLER_0_160_1173 ();
 sg13g2_fill_8 FILLER_0_160_1183 ();
 sg13g2_fill_8 FILLER_0_160_1191 ();
 sg13g2_fill_1 FILLER_0_160_1199 ();
 sg13g2_fill_2 FILLER_0_160_1221 ();
 sg13g2_fill_2 FILLER_0_160_1227 ();
 sg13g2_fill_4 FILLER_0_160_1234 ();
 sg13g2_fill_1 FILLER_0_160_1238 ();
 sg13g2_fill_8 FILLER_0_160_1243 ();
 sg13g2_fill_8 FILLER_0_160_1251 ();
 sg13g2_fill_8 FILLER_0_160_1259 ();
 sg13g2_fill_8 FILLER_0_160_1267 ();
 sg13g2_fill_8 FILLER_0_160_1275 ();
 sg13g2_fill_8 FILLER_0_160_1283 ();
 sg13g2_fill_4 FILLER_0_160_1291 ();
 sg13g2_fill_2 FILLER_0_160_1295 ();
 sg13g2_fill_8 FILLER_0_161_0 ();
 sg13g2_fill_8 FILLER_0_161_8 ();
 sg13g2_fill_8 FILLER_0_161_16 ();
 sg13g2_fill_8 FILLER_0_161_24 ();
 sg13g2_fill_8 FILLER_0_161_32 ();
 sg13g2_fill_8 FILLER_0_161_40 ();
 sg13g2_fill_8 FILLER_0_161_48 ();
 sg13g2_fill_8 FILLER_0_161_56 ();
 sg13g2_fill_8 FILLER_0_161_64 ();
 sg13g2_fill_8 FILLER_0_161_72 ();
 sg13g2_fill_8 FILLER_0_161_80 ();
 sg13g2_fill_8 FILLER_0_161_88 ();
 sg13g2_fill_8 FILLER_0_161_96 ();
 sg13g2_fill_8 FILLER_0_161_104 ();
 sg13g2_fill_8 FILLER_0_161_112 ();
 sg13g2_fill_8 FILLER_0_161_120 ();
 sg13g2_fill_8 FILLER_0_161_128 ();
 sg13g2_fill_8 FILLER_0_161_136 ();
 sg13g2_fill_8 FILLER_0_161_144 ();
 sg13g2_fill_8 FILLER_0_161_152 ();
 sg13g2_fill_8 FILLER_0_161_160 ();
 sg13g2_fill_8 FILLER_0_161_168 ();
 sg13g2_fill_8 FILLER_0_161_176 ();
 sg13g2_fill_8 FILLER_0_161_184 ();
 sg13g2_fill_8 FILLER_0_161_192 ();
 sg13g2_fill_8 FILLER_0_161_200 ();
 sg13g2_fill_8 FILLER_0_161_208 ();
 sg13g2_fill_8 FILLER_0_161_216 ();
 sg13g2_fill_8 FILLER_0_161_224 ();
 sg13g2_fill_8 FILLER_0_161_232 ();
 sg13g2_fill_8 FILLER_0_161_240 ();
 sg13g2_fill_8 FILLER_0_161_248 ();
 sg13g2_fill_8 FILLER_0_161_256 ();
 sg13g2_fill_8 FILLER_0_161_264 ();
 sg13g2_fill_8 FILLER_0_161_272 ();
 sg13g2_fill_8 FILLER_0_161_280 ();
 sg13g2_fill_8 FILLER_0_161_288 ();
 sg13g2_fill_8 FILLER_0_161_296 ();
 sg13g2_fill_8 FILLER_0_161_304 ();
 sg13g2_fill_8 FILLER_0_161_312 ();
 sg13g2_fill_8 FILLER_0_161_320 ();
 sg13g2_fill_8 FILLER_0_161_328 ();
 sg13g2_fill_8 FILLER_0_161_336 ();
 sg13g2_fill_8 FILLER_0_161_344 ();
 sg13g2_fill_8 FILLER_0_161_352 ();
 sg13g2_fill_8 FILLER_0_161_360 ();
 sg13g2_fill_8 FILLER_0_161_368 ();
 sg13g2_fill_8 FILLER_0_161_376 ();
 sg13g2_fill_8 FILLER_0_161_384 ();
 sg13g2_fill_8 FILLER_0_161_392 ();
 sg13g2_fill_8 FILLER_0_161_400 ();
 sg13g2_fill_8 FILLER_0_161_408 ();
 sg13g2_fill_8 FILLER_0_161_416 ();
 sg13g2_fill_8 FILLER_0_161_424 ();
 sg13g2_fill_8 FILLER_0_161_432 ();
 sg13g2_fill_8 FILLER_0_161_440 ();
 sg13g2_fill_8 FILLER_0_161_448 ();
 sg13g2_fill_8 FILLER_0_161_456 ();
 sg13g2_fill_8 FILLER_0_161_464 ();
 sg13g2_fill_8 FILLER_0_161_472 ();
 sg13g2_fill_8 FILLER_0_161_480 ();
 sg13g2_fill_8 FILLER_0_161_488 ();
 sg13g2_fill_8 FILLER_0_161_496 ();
 sg13g2_fill_8 FILLER_0_161_504 ();
 sg13g2_fill_8 FILLER_0_161_512 ();
 sg13g2_fill_8 FILLER_0_161_520 ();
 sg13g2_fill_8 FILLER_0_161_528 ();
 sg13g2_fill_8 FILLER_0_161_536 ();
 sg13g2_fill_8 FILLER_0_161_544 ();
 sg13g2_fill_8 FILLER_0_161_552 ();
 sg13g2_fill_8 FILLER_0_161_560 ();
 sg13g2_fill_2 FILLER_0_161_572 ();
 sg13g2_fill_2 FILLER_0_161_579 ();
 sg13g2_fill_8 FILLER_0_161_607 ();
 sg13g2_fill_8 FILLER_0_161_615 ();
 sg13g2_fill_8 FILLER_0_161_623 ();
 sg13g2_fill_8 FILLER_0_161_631 ();
 sg13g2_fill_4 FILLER_0_161_639 ();
 sg13g2_fill_2 FILLER_0_161_648 ();
 sg13g2_fill_2 FILLER_0_161_676 ();
 sg13g2_fill_2 FILLER_0_161_683 ();
 sg13g2_fill_2 FILLER_0_161_693 ();
 sg13g2_fill_1 FILLER_0_161_695 ();
 sg13g2_fill_4 FILLER_0_161_700 ();
 sg13g2_fill_2 FILLER_0_161_704 ();
 sg13g2_fill_1 FILLER_0_161_706 ();
 sg13g2_fill_4 FILLER_0_161_733 ();
 sg13g2_fill_2 FILLER_0_161_737 ();
 sg13g2_fill_1 FILLER_0_161_739 ();
 sg13g2_fill_2 FILLER_0_161_745 ();
 sg13g2_fill_2 FILLER_0_161_751 ();
 sg13g2_fill_1 FILLER_0_161_753 ();
 sg13g2_fill_2 FILLER_0_161_759 ();
 sg13g2_fill_1 FILLER_0_161_761 ();
 sg13g2_fill_2 FILLER_0_161_766 ();
 sg13g2_fill_1 FILLER_0_161_768 ();
 sg13g2_fill_2 FILLER_0_161_774 ();
 sg13g2_fill_1 FILLER_0_161_776 ();
 sg13g2_fill_4 FILLER_0_161_781 ();
 sg13g2_fill_1 FILLER_0_161_785 ();
 sg13g2_fill_8 FILLER_0_161_791 ();
 sg13g2_fill_8 FILLER_0_161_804 ();
 sg13g2_fill_4 FILLER_0_161_817 ();
 sg13g2_fill_2 FILLER_0_161_821 ();
 sg13g2_fill_1 FILLER_0_161_823 ();
 sg13g2_fill_4 FILLER_0_161_829 ();
 sg13g2_fill_1 FILLER_0_161_833 ();
 sg13g2_fill_4 FILLER_0_161_838 ();
 sg13g2_fill_2 FILLER_0_161_842 ();
 sg13g2_fill_1 FILLER_0_161_844 ();
 sg13g2_fill_2 FILLER_0_161_850 ();
 sg13g2_fill_1 FILLER_0_161_852 ();
 sg13g2_fill_4 FILLER_0_161_861 ();
 sg13g2_fill_8 FILLER_0_161_873 ();
 sg13g2_fill_2 FILLER_0_161_881 ();
 sg13g2_fill_1 FILLER_0_161_883 ();
 sg13g2_fill_2 FILLER_0_161_892 ();
 sg13g2_fill_2 FILLER_0_161_899 ();
 sg13g2_fill_2 FILLER_0_161_927 ();
 sg13g2_fill_2 FILLER_0_161_933 ();
 sg13g2_fill_2 FILLER_0_161_945 ();
 sg13g2_fill_1 FILLER_0_161_947 ();
 sg13g2_fill_2 FILLER_0_161_952 ();
 sg13g2_fill_2 FILLER_0_161_959 ();
 sg13g2_fill_8 FILLER_0_161_966 ();
 sg13g2_fill_2 FILLER_0_161_974 ();
 sg13g2_fill_4 FILLER_0_161_980 ();
 sg13g2_fill_4 FILLER_0_161_1010 ();
 sg13g2_fill_2 FILLER_0_161_1014 ();
 sg13g2_fill_4 FILLER_0_161_1021 ();
 sg13g2_fill_2 FILLER_0_161_1025 ();
 sg13g2_fill_4 FILLER_0_161_1053 ();
 sg13g2_fill_1 FILLER_0_161_1057 ();
 sg13g2_fill_2 FILLER_0_161_1063 ();
 sg13g2_fill_4 FILLER_0_161_1091 ();
 sg13g2_fill_1 FILLER_0_161_1095 ();
 sg13g2_fill_4 FILLER_0_161_1122 ();
 sg13g2_fill_1 FILLER_0_161_1126 ();
 sg13g2_fill_8 FILLER_0_161_1132 ();
 sg13g2_fill_4 FILLER_0_161_1140 ();
 sg13g2_fill_4 FILLER_0_161_1149 ();
 sg13g2_fill_2 FILLER_0_161_1153 ();
 sg13g2_fill_4 FILLER_0_161_1159 ();
 sg13g2_fill_2 FILLER_0_161_1163 ();
 sg13g2_fill_4 FILLER_0_161_1186 ();
 sg13g2_fill_2 FILLER_0_161_1190 ();
 sg13g2_fill_2 FILLER_0_161_1197 ();
 sg13g2_fill_8 FILLER_0_161_1203 ();
 sg13g2_fill_8 FILLER_0_161_1211 ();
 sg13g2_fill_8 FILLER_0_161_1219 ();
 sg13g2_fill_2 FILLER_0_161_1227 ();
 sg13g2_fill_8 FILLER_0_161_1255 ();
 sg13g2_fill_8 FILLER_0_161_1263 ();
 sg13g2_fill_8 FILLER_0_161_1271 ();
 sg13g2_fill_8 FILLER_0_161_1279 ();
 sg13g2_fill_8 FILLER_0_161_1287 ();
 sg13g2_fill_2 FILLER_0_161_1295 ();
 sg13g2_fill_8 FILLER_0_162_0 ();
 sg13g2_fill_8 FILLER_0_162_8 ();
 sg13g2_fill_8 FILLER_0_162_16 ();
 sg13g2_fill_8 FILLER_0_162_24 ();
 sg13g2_fill_8 FILLER_0_162_32 ();
 sg13g2_fill_8 FILLER_0_162_40 ();
 sg13g2_fill_8 FILLER_0_162_48 ();
 sg13g2_fill_8 FILLER_0_162_56 ();
 sg13g2_fill_8 FILLER_0_162_64 ();
 sg13g2_fill_8 FILLER_0_162_72 ();
 sg13g2_fill_8 FILLER_0_162_80 ();
 sg13g2_fill_8 FILLER_0_162_88 ();
 sg13g2_fill_8 FILLER_0_162_96 ();
 sg13g2_fill_8 FILLER_0_162_104 ();
 sg13g2_fill_8 FILLER_0_162_112 ();
 sg13g2_fill_8 FILLER_0_162_120 ();
 sg13g2_fill_8 FILLER_0_162_128 ();
 sg13g2_fill_8 FILLER_0_162_136 ();
 sg13g2_fill_8 FILLER_0_162_144 ();
 sg13g2_fill_8 FILLER_0_162_152 ();
 sg13g2_fill_8 FILLER_0_162_160 ();
 sg13g2_fill_8 FILLER_0_162_168 ();
 sg13g2_fill_8 FILLER_0_162_176 ();
 sg13g2_fill_8 FILLER_0_162_184 ();
 sg13g2_fill_8 FILLER_0_162_192 ();
 sg13g2_fill_8 FILLER_0_162_200 ();
 sg13g2_fill_8 FILLER_0_162_208 ();
 sg13g2_fill_8 FILLER_0_162_216 ();
 sg13g2_fill_8 FILLER_0_162_224 ();
 sg13g2_fill_8 FILLER_0_162_232 ();
 sg13g2_fill_8 FILLER_0_162_240 ();
 sg13g2_fill_8 FILLER_0_162_248 ();
 sg13g2_fill_8 FILLER_0_162_256 ();
 sg13g2_fill_8 FILLER_0_162_264 ();
 sg13g2_fill_8 FILLER_0_162_272 ();
 sg13g2_fill_8 FILLER_0_162_280 ();
 sg13g2_fill_8 FILLER_0_162_288 ();
 sg13g2_fill_8 FILLER_0_162_296 ();
 sg13g2_fill_8 FILLER_0_162_304 ();
 sg13g2_fill_8 FILLER_0_162_312 ();
 sg13g2_fill_8 FILLER_0_162_320 ();
 sg13g2_fill_8 FILLER_0_162_328 ();
 sg13g2_fill_8 FILLER_0_162_336 ();
 sg13g2_fill_8 FILLER_0_162_344 ();
 sg13g2_fill_8 FILLER_0_162_352 ();
 sg13g2_fill_8 FILLER_0_162_360 ();
 sg13g2_fill_8 FILLER_0_162_368 ();
 sg13g2_fill_8 FILLER_0_162_376 ();
 sg13g2_fill_8 FILLER_0_162_384 ();
 sg13g2_fill_8 FILLER_0_162_392 ();
 sg13g2_fill_8 FILLER_0_162_400 ();
 sg13g2_fill_8 FILLER_0_162_408 ();
 sg13g2_fill_8 FILLER_0_162_416 ();
 sg13g2_fill_8 FILLER_0_162_424 ();
 sg13g2_fill_8 FILLER_0_162_432 ();
 sg13g2_fill_8 FILLER_0_162_440 ();
 sg13g2_fill_8 FILLER_0_162_448 ();
 sg13g2_fill_8 FILLER_0_162_456 ();
 sg13g2_fill_8 FILLER_0_162_464 ();
 sg13g2_fill_8 FILLER_0_162_472 ();
 sg13g2_fill_8 FILLER_0_162_480 ();
 sg13g2_fill_8 FILLER_0_162_488 ();
 sg13g2_fill_8 FILLER_0_162_496 ();
 sg13g2_fill_8 FILLER_0_162_504 ();
 sg13g2_fill_8 FILLER_0_162_512 ();
 sg13g2_fill_8 FILLER_0_162_520 ();
 sg13g2_fill_8 FILLER_0_162_528 ();
 sg13g2_fill_8 FILLER_0_162_536 ();
 sg13g2_fill_8 FILLER_0_162_544 ();
 sg13g2_fill_8 FILLER_0_162_552 ();
 sg13g2_fill_8 FILLER_0_162_560 ();
 sg13g2_fill_8 FILLER_0_162_568 ();
 sg13g2_fill_8 FILLER_0_162_576 ();
 sg13g2_fill_8 FILLER_0_162_584 ();
 sg13g2_fill_8 FILLER_0_162_592 ();
 sg13g2_fill_8 FILLER_0_162_600 ();
 sg13g2_fill_8 FILLER_0_162_608 ();
 sg13g2_fill_8 FILLER_0_162_616 ();
 sg13g2_fill_8 FILLER_0_162_624 ();
 sg13g2_fill_2 FILLER_0_162_632 ();
 sg13g2_fill_1 FILLER_0_162_634 ();
 sg13g2_fill_8 FILLER_0_162_661 ();
 sg13g2_fill_8 FILLER_0_162_669 ();
 sg13g2_fill_8 FILLER_0_162_677 ();
 sg13g2_fill_4 FILLER_0_162_685 ();
 sg13g2_fill_2 FILLER_0_162_689 ();
 sg13g2_fill_4 FILLER_0_162_696 ();
 sg13g2_fill_2 FILLER_0_162_700 ();
 sg13g2_fill_1 FILLER_0_162_702 ();
 sg13g2_fill_2 FILLER_0_162_708 ();
 sg13g2_fill_8 FILLER_0_162_715 ();
 sg13g2_fill_4 FILLER_0_162_723 ();
 sg13g2_fill_2 FILLER_0_162_727 ();
 sg13g2_fill_8 FILLER_0_162_733 ();
 sg13g2_fill_4 FILLER_0_162_741 ();
 sg13g2_fill_1 FILLER_0_162_745 ();
 sg13g2_fill_4 FILLER_0_162_772 ();
 sg13g2_fill_2 FILLER_0_162_776 ();
 sg13g2_fill_2 FILLER_0_162_783 ();
 sg13g2_fill_1 FILLER_0_162_785 ();
 sg13g2_fill_8 FILLER_0_162_812 ();
 sg13g2_fill_4 FILLER_0_162_820 ();
 sg13g2_fill_1 FILLER_0_162_824 ();
 sg13g2_fill_4 FILLER_0_162_851 ();
 sg13g2_fill_1 FILLER_0_162_855 ();
 sg13g2_fill_4 FILLER_0_162_882 ();
 sg13g2_fill_1 FILLER_0_162_886 ();
 sg13g2_fill_2 FILLER_0_162_892 ();
 sg13g2_fill_2 FILLER_0_162_899 ();
 sg13g2_fill_4 FILLER_0_162_906 ();
 sg13g2_fill_1 FILLER_0_162_910 ();
 sg13g2_fill_4 FILLER_0_162_915 ();
 sg13g2_fill_2 FILLER_0_162_924 ();
 sg13g2_fill_1 FILLER_0_162_926 ();
 sg13g2_fill_2 FILLER_0_162_931 ();
 sg13g2_fill_2 FILLER_0_162_937 ();
 sg13g2_fill_2 FILLER_0_162_943 ();
 sg13g2_fill_8 FILLER_0_162_949 ();
 sg13g2_fill_8 FILLER_0_162_957 ();
 sg13g2_fill_8 FILLER_0_162_965 ();
 sg13g2_fill_4 FILLER_0_162_973 ();
 sg13g2_fill_2 FILLER_0_162_977 ();
 sg13g2_fill_8 FILLER_0_162_1000 ();
 sg13g2_fill_2 FILLER_0_162_1034 ();
 sg13g2_fill_4 FILLER_0_162_1041 ();
 sg13g2_fill_1 FILLER_0_162_1045 ();
 sg13g2_fill_8 FILLER_0_162_1050 ();
 sg13g2_fill_4 FILLER_0_162_1058 ();
 sg13g2_fill_2 FILLER_0_162_1067 ();
 sg13g2_fill_8 FILLER_0_162_1073 ();
 sg13g2_fill_8 FILLER_0_162_1087 ();
 sg13g2_fill_4 FILLER_0_162_1095 ();
 sg13g2_fill_2 FILLER_0_162_1104 ();
 sg13g2_fill_1 FILLER_0_162_1106 ();
 sg13g2_fill_8 FILLER_0_162_1111 ();
 sg13g2_fill_4 FILLER_0_162_1119 ();
 sg13g2_fill_2 FILLER_0_162_1123 ();
 sg13g2_fill_8 FILLER_0_162_1130 ();
 sg13g2_fill_8 FILLER_0_162_1138 ();
 sg13g2_fill_2 FILLER_0_162_1146 ();
 sg13g2_fill_2 FILLER_0_162_1174 ();
 sg13g2_fill_4 FILLER_0_162_1181 ();
 sg13g2_fill_8 FILLER_0_162_1211 ();
 sg13g2_fill_8 FILLER_0_162_1219 ();
 sg13g2_fill_8 FILLER_0_162_1227 ();
 sg13g2_fill_8 FILLER_0_162_1235 ();
 sg13g2_fill_8 FILLER_0_162_1243 ();
 sg13g2_fill_8 FILLER_0_162_1251 ();
 sg13g2_fill_8 FILLER_0_162_1259 ();
 sg13g2_fill_8 FILLER_0_162_1267 ();
 sg13g2_fill_8 FILLER_0_162_1275 ();
 sg13g2_fill_8 FILLER_0_162_1283 ();
 sg13g2_fill_4 FILLER_0_162_1291 ();
 sg13g2_fill_2 FILLER_0_162_1295 ();
 sg13g2_fill_8 FILLER_0_163_0 ();
 sg13g2_fill_8 FILLER_0_163_8 ();
 sg13g2_fill_8 FILLER_0_163_16 ();
 sg13g2_fill_8 FILLER_0_163_24 ();
 sg13g2_fill_8 FILLER_0_163_32 ();
 sg13g2_fill_8 FILLER_0_163_40 ();
 sg13g2_fill_8 FILLER_0_163_48 ();
 sg13g2_fill_8 FILLER_0_163_56 ();
 sg13g2_fill_8 FILLER_0_163_64 ();
 sg13g2_fill_8 FILLER_0_163_72 ();
 sg13g2_fill_8 FILLER_0_163_80 ();
 sg13g2_fill_8 FILLER_0_163_88 ();
 sg13g2_fill_8 FILLER_0_163_96 ();
 sg13g2_fill_8 FILLER_0_163_104 ();
 sg13g2_fill_8 FILLER_0_163_112 ();
 sg13g2_fill_8 FILLER_0_163_120 ();
 sg13g2_fill_8 FILLER_0_163_128 ();
 sg13g2_fill_8 FILLER_0_163_136 ();
 sg13g2_fill_8 FILLER_0_163_144 ();
 sg13g2_fill_8 FILLER_0_163_152 ();
 sg13g2_fill_8 FILLER_0_163_160 ();
 sg13g2_fill_8 FILLER_0_163_168 ();
 sg13g2_fill_8 FILLER_0_163_176 ();
 sg13g2_fill_8 FILLER_0_163_184 ();
 sg13g2_fill_8 FILLER_0_163_192 ();
 sg13g2_fill_8 FILLER_0_163_200 ();
 sg13g2_fill_8 FILLER_0_163_208 ();
 sg13g2_fill_8 FILLER_0_163_216 ();
 sg13g2_fill_8 FILLER_0_163_224 ();
 sg13g2_fill_8 FILLER_0_163_232 ();
 sg13g2_fill_8 FILLER_0_163_240 ();
 sg13g2_fill_8 FILLER_0_163_248 ();
 sg13g2_fill_8 FILLER_0_163_256 ();
 sg13g2_fill_8 FILLER_0_163_264 ();
 sg13g2_fill_8 FILLER_0_163_272 ();
 sg13g2_fill_8 FILLER_0_163_280 ();
 sg13g2_fill_8 FILLER_0_163_288 ();
 sg13g2_fill_8 FILLER_0_163_296 ();
 sg13g2_fill_8 FILLER_0_163_304 ();
 sg13g2_fill_8 FILLER_0_163_312 ();
 sg13g2_fill_8 FILLER_0_163_320 ();
 sg13g2_fill_8 FILLER_0_163_328 ();
 sg13g2_fill_8 FILLER_0_163_336 ();
 sg13g2_fill_8 FILLER_0_163_344 ();
 sg13g2_fill_8 FILLER_0_163_352 ();
 sg13g2_fill_8 FILLER_0_163_360 ();
 sg13g2_fill_8 FILLER_0_163_368 ();
 sg13g2_fill_8 FILLER_0_163_376 ();
 sg13g2_fill_8 FILLER_0_163_384 ();
 sg13g2_fill_8 FILLER_0_163_392 ();
 sg13g2_fill_8 FILLER_0_163_400 ();
 sg13g2_fill_8 FILLER_0_163_408 ();
 sg13g2_fill_8 FILLER_0_163_416 ();
 sg13g2_fill_8 FILLER_0_163_424 ();
 sg13g2_fill_8 FILLER_0_163_432 ();
 sg13g2_fill_8 FILLER_0_163_440 ();
 sg13g2_fill_8 FILLER_0_163_448 ();
 sg13g2_fill_8 FILLER_0_163_456 ();
 sg13g2_fill_8 FILLER_0_163_464 ();
 sg13g2_fill_8 FILLER_0_163_472 ();
 sg13g2_fill_8 FILLER_0_163_480 ();
 sg13g2_fill_8 FILLER_0_163_488 ();
 sg13g2_fill_8 FILLER_0_163_496 ();
 sg13g2_fill_8 FILLER_0_163_504 ();
 sg13g2_fill_8 FILLER_0_163_512 ();
 sg13g2_fill_8 FILLER_0_163_520 ();
 sg13g2_fill_8 FILLER_0_163_528 ();
 sg13g2_fill_8 FILLER_0_163_536 ();
 sg13g2_fill_4 FILLER_0_163_544 ();
 sg13g2_fill_2 FILLER_0_163_548 ();
 sg13g2_fill_1 FILLER_0_163_550 ();
 sg13g2_fill_8 FILLER_0_163_555 ();
 sg13g2_fill_8 FILLER_0_163_563 ();
 sg13g2_fill_8 FILLER_0_163_571 ();
 sg13g2_fill_8 FILLER_0_163_579 ();
 sg13g2_fill_8 FILLER_0_163_587 ();
 sg13g2_fill_8 FILLER_0_163_595 ();
 sg13g2_fill_8 FILLER_0_163_603 ();
 sg13g2_fill_8 FILLER_0_163_611 ();
 sg13g2_fill_8 FILLER_0_163_619 ();
 sg13g2_fill_8 FILLER_0_163_627 ();
 sg13g2_fill_2 FILLER_0_163_635 ();
 sg13g2_fill_2 FILLER_0_163_642 ();
 sg13g2_fill_8 FILLER_0_163_648 ();
 sg13g2_fill_8 FILLER_0_163_656 ();
 sg13g2_fill_8 FILLER_0_163_664 ();
 sg13g2_fill_8 FILLER_0_163_672 ();
 sg13g2_fill_8 FILLER_0_163_680 ();
 sg13g2_fill_8 FILLER_0_163_688 ();
 sg13g2_fill_8 FILLER_0_163_696 ();
 sg13g2_fill_8 FILLER_0_163_704 ();
 sg13g2_fill_8 FILLER_0_163_712 ();
 sg13g2_fill_8 FILLER_0_163_720 ();
 sg13g2_fill_8 FILLER_0_163_728 ();
 sg13g2_fill_8 FILLER_0_163_736 ();
 sg13g2_fill_8 FILLER_0_163_744 ();
 sg13g2_fill_8 FILLER_0_163_752 ();
 sg13g2_fill_8 FILLER_0_163_760 ();
 sg13g2_fill_8 FILLER_0_163_768 ();
 sg13g2_fill_8 FILLER_0_163_776 ();
 sg13g2_fill_2 FILLER_0_163_784 ();
 sg13g2_fill_4 FILLER_0_163_790 ();
 sg13g2_fill_2 FILLER_0_163_794 ();
 sg13g2_fill_1 FILLER_0_163_796 ();
 sg13g2_fill_4 FILLER_0_163_801 ();
 sg13g2_fill_8 FILLER_0_163_809 ();
 sg13g2_fill_8 FILLER_0_163_817 ();
 sg13g2_fill_8 FILLER_0_163_825 ();
 sg13g2_fill_4 FILLER_0_163_833 ();
 sg13g2_fill_1 FILLER_0_163_837 ();
 sg13g2_fill_8 FILLER_0_163_843 ();
 sg13g2_fill_4 FILLER_0_163_851 ();
 sg13g2_fill_2 FILLER_0_163_860 ();
 sg13g2_fill_2 FILLER_0_163_866 ();
 sg13g2_fill_2 FILLER_0_163_873 ();
 sg13g2_fill_2 FILLER_0_163_879 ();
 sg13g2_fill_2 FILLER_0_163_885 ();
 sg13g2_fill_1 FILLER_0_163_887 ();
 sg13g2_fill_2 FILLER_0_163_892 ();
 sg13g2_fill_2 FILLER_0_163_898 ();
 sg13g2_fill_2 FILLER_0_163_904 ();
 sg13g2_fill_2 FILLER_0_163_910 ();
 sg13g2_fill_2 FILLER_0_163_917 ();
 sg13g2_fill_2 FILLER_0_163_923 ();
 sg13g2_fill_2 FILLER_0_163_930 ();
 sg13g2_fill_8 FILLER_0_163_936 ();
 sg13g2_fill_2 FILLER_0_163_944 ();
 sg13g2_fill_8 FILLER_0_163_950 ();
 sg13g2_fill_8 FILLER_0_163_958 ();
 sg13g2_fill_8 FILLER_0_163_966 ();
 sg13g2_fill_8 FILLER_0_163_974 ();
 sg13g2_fill_8 FILLER_0_163_982 ();
 sg13g2_fill_8 FILLER_0_163_990 ();
 sg13g2_fill_8 FILLER_0_163_998 ();
 sg13g2_fill_4 FILLER_0_163_1006 ();
 sg13g2_fill_8 FILLER_0_163_1015 ();
 sg13g2_fill_8 FILLER_0_163_1023 ();
 sg13g2_fill_8 FILLER_0_163_1031 ();
 sg13g2_fill_8 FILLER_0_163_1039 ();
 sg13g2_fill_8 FILLER_0_163_1047 ();
 sg13g2_fill_8 FILLER_0_163_1055 ();
 sg13g2_fill_8 FILLER_0_163_1063 ();
 sg13g2_fill_8 FILLER_0_163_1071 ();
 sg13g2_fill_8 FILLER_0_163_1079 ();
 sg13g2_fill_8 FILLER_0_163_1087 ();
 sg13g2_fill_8 FILLER_0_163_1095 ();
 sg13g2_fill_8 FILLER_0_163_1103 ();
 sg13g2_fill_8 FILLER_0_163_1111 ();
 sg13g2_fill_8 FILLER_0_163_1119 ();
 sg13g2_fill_8 FILLER_0_163_1127 ();
 sg13g2_fill_8 FILLER_0_163_1135 ();
 sg13g2_fill_8 FILLER_0_163_1143 ();
 sg13g2_fill_8 FILLER_0_163_1151 ();
 sg13g2_fill_8 FILLER_0_163_1159 ();
 sg13g2_fill_1 FILLER_0_163_1167 ();
 sg13g2_fill_8 FILLER_0_163_1172 ();
 sg13g2_fill_8 FILLER_0_163_1180 ();
 sg13g2_fill_8 FILLER_0_163_1188 ();
 sg13g2_fill_8 FILLER_0_163_1196 ();
 sg13g2_fill_8 FILLER_0_163_1204 ();
 sg13g2_fill_8 FILLER_0_163_1212 ();
 sg13g2_fill_8 FILLER_0_163_1220 ();
 sg13g2_fill_8 FILLER_0_163_1228 ();
 sg13g2_fill_8 FILLER_0_163_1236 ();
 sg13g2_fill_8 FILLER_0_163_1244 ();
 sg13g2_fill_8 FILLER_0_163_1252 ();
 sg13g2_fill_8 FILLER_0_163_1260 ();
 sg13g2_fill_8 FILLER_0_163_1268 ();
 sg13g2_fill_8 FILLER_0_163_1276 ();
 sg13g2_fill_8 FILLER_0_163_1284 ();
 sg13g2_fill_4 FILLER_0_163_1292 ();
 sg13g2_fill_1 FILLER_0_163_1296 ();
endmodule
