** sch_path: /home/ac3e/Documents/ihp_design/klayout/netlist/rdiv.sch
.subckt rdiv vout vss in_p
*.PININFO vout:B vss:B in_p:B
R2 vss in_p rhigh w=0.5e-6 l=30e-6 m=1 b=0
R1 in_p vout rhigh w=0.5e-6 l=10e-6 m=1 b=0
.ends
.end
