** sch_path: /home/ac3e/Documents/ihp_design/klayout/netlist/OTA_without_rcomp.sch
.subckt OTA iref vin_n vin_p vdd vss vout
*.PININFO iref:I vin_n:I vin_p:I vdd:B vss:B vout:O
M1 net1 vin_n net2 1 sg13_lv_nmos W=15u L=2u ng=1 m=1
M2 net3 vin_p net2 1 sg13_lv_nmos W=15u L=2u ng=1 m=1
M3 net3 net1 vdd 2 sg13_lv_pmos W=2u L=1u ng=1 m=1
M4 net1 net1 vdd 2 sg13_lv_pmos W=2u L=1u ng=1 m=1
M5 net2 iref vss 1 sg13_lv_nmos W=6u L=2u ng=1 m=1
M8 iref iref vss 1 sg13_lv_nmos W=6u L=2u ng=1 m=1
M6 vout net3 vdd 2 sg13_lv_pmos W=20u L=0.5u ng=1 m=1
M7 vout iref vss 1 sg13_lv_nmos W=24u L=2u ng=1 m=1
C2 vout net4 cap_cmim W=45.0e-6 L=45.0e-6 MF=1
R2 net3 net4 rhigh w=0.5e-6 l=3.5e-6 m=1 b=0
.ends
.end
