** sch_path: /home/herman/github/KrzysztofHerman/IHP-Open-DesignLib/ts_pr_May2024/design_data/xschem/transmission_gate_tb.sch
.subckt transmission_gate_tb

Vpow net1 GND 1.2
Vp net1 net2 0
.save i(vp)
Vin V_in GND dc=0 ac=1 sin(0, 200m, 20meg, 0, 0)
Ven en_in GND pulse(0 1.2 0 1p 1p 50n 100n)
C1 V_out GND 10p m=1
x1 net2 V_in V_out GND en_in tgate
**** begin user architecture code

.lib /home/herman/github/KrzysztofHerman/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /home/herman/github/KrzysztofHerman/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.include /home/herman/github/KrzysztofHerman/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/diodes.lib
.include /home/herman/github/KrzysztofHerman/IHP-Open-PDK/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27
.control
pre_osdi ./psp103_nqs.osdi
save all
tran 100p 120n
write tran_res_temp.raw
.endc


**** end user architecture code
.ends

* expanding   symbol:  tgate.sym # of pins=5
** sym_path: /home/herman/github/KrzysztofHerman/IHP-Open-DesignLib/ts_pr_May2024/design_data/xschem/tgate.sym
** sch_path: /home/herman/github/KrzysztofHerman/IHP-Open-DesignLib/ts_pr_May2024/design_data/xschem/tgate.sch
.subckt tgate vdd inout_1 inout_2 vss en
*.PININFO inout_1:B inout_2:B en:I vdd:B vss:B
M1 inout_2 net1 inout_1 sub sg13_lv_nmos L=0.130u W=5.0u ng=5 m=1
M2 inout_1 en inout_2 nwell sg13_lv_pmos L=0.130u W=5.0u ng=5 m=1
R1 vss sub ptap1 l=780n w=780n
R2 vdd nwell ntap1 l=780n w=780n
M3 net1 en vss sub sg13_lv_nmos L=0.130u W=0.740u ng=1 m=1
M4 net1 en vdd nwell sg13_lv_pmos L=0.130u W=1.120u ng=1 m=1
D1 sub en dantenna l=780n w=780n
D2 en nwell dpantenna l=780n w=780n
.ends

.GLOBAL GND
.end
